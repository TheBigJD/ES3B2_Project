
//////////////////////////////////////////////////////////////////////////////////
//Solid_block
//////////////////////////////////////////////////////////////////////////////////


module Pacman(

  input Master_Clock_In,
  input [9 : 0] xInput,
  input [9 : 0] yInput,
  output reg [11:0] ColourData = 12'h000

);

(* rom_style = "block" *)

reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

always @(posedge Master_Clock_In)
begin
  a = xInput % 32;
  b = yInput % 32;

Inputs = {a, b};

    case(Inputs)
    
20'b00000000000000000000 : ColourData = 12'hFFF;
20'b00000000010000000000 : ColourData = 12'hFFF;
20'b00000000100000000000 : ColourData = 12'hFFF;
20'b00000000110000000000 : ColourData = 12'hFFF;
20'b00000001000000000000 : ColourData = 12'hFFF;
20'b00000001010000000000 : ColourData = 12'hFFF;
20'b00000001100000000000 : ColourData = 12'hFFF;
20'b00000001110000000000 : ColourData = 12'hFFF;
20'b00000010000000000000 : ColourData = 12'hFFF;
20'b00000010010000000000 : ColourData = 12'hFFF;
20'b00000010100000000000 : ColourData = 12'hFFF;
20'b00000010110000000000 : ColourData = 12'hFFF;
20'b00000011000000000000 : ColourData = 12'hFFF;
20'b00000011010000000000 : ColourData = 12'hFFF;
20'b00000011100000000000 : ColourData = 12'hFFF;
20'b00000011110000000000 : ColourData = 12'hFFF;
20'b00000100000000000000 : ColourData = 12'hFFF;
20'b00000100010000000000 : ColourData = 12'hFFF;
20'b00000100100000000000 : ColourData = 12'hFFF;
20'b00000100110000000000 : ColourData = 12'hFFF;
20'b00000101000000000000 : ColourData = 12'hFFF;
20'b00000101010000000000 : ColourData = 12'hFFF;
20'b00000101100000000000 : ColourData = 12'hFFF;
20'b00000101110000000000 : ColourData = 12'hFFF;
20'b00000110000000000000 : ColourData = 12'hFFF;
20'b00000000000000000001 : ColourData = 12'hFFF;
20'b00000000010000000001 : ColourData = 12'hFFF;
20'b00000000100000000001 : ColourData = 12'hFFF;
20'b00000000110000000001 : ColourData = 12'hFFF;
20'b00000001000000000001 : ColourData = 12'hFFF;
20'b00000001010000000001 : ColourData = 12'hFFF;
20'b00000001100000000001 : ColourData = 12'hFFF;
20'b00000001110000000001 : ColourData = 12'hFFF;
20'b00000010000000000001 : ColourData = 12'hFFF;
20'b00000010010000000001 : ColourData = 12'hDF0;
20'b00000010100000000001 : ColourData = 12'hDF0;
20'b00000010110000000001 : ColourData = 12'hDF0;
20'b00000011000000000001 : ColourData = 12'hDF0;
20'b00000011010000000001 : ColourData = 12'hDF0;
20'b00000011100000000001 : ColourData = 12'hDF0;
20'b00000011110000000001 : ColourData = 12'hDF0;
20'b00000100000000000001 : ColourData = 12'hFFF;
20'b00000100010000000001 : ColourData = 12'hFFF;
20'b00000100100000000001 : ColourData = 12'hFFF;
20'b00000100110000000001 : ColourData = 12'hFFF;
20'b00000101000000000001 : ColourData = 12'hFFF;
20'b00000101010000000001 : ColourData = 12'hFFF;
20'b00000101100000000001 : ColourData = 12'hFFF;
20'b00000101110000000001 : ColourData = 12'hFFF;
20'b00000110000000000001 : ColourData = 12'hFFF;
20'b00000000000000000010 : ColourData = 12'hFFF;
20'b00000000010000000010 : ColourData = 12'hFFF;
20'b00000000100000000010 : ColourData = 12'hFFF;
20'b00000000110000000010 : ColourData = 12'hFFF;
20'b00000001000000000010 : ColourData = 12'hFFF;
20'b00000001010000000010 : ColourData = 12'hFFF;
20'b00000001100000000010 : ColourData = 12'hFFF;
20'b00000001110000000010 : ColourData = 12'hDF0;
20'b00000010000000000010 : ColourData = 12'hDF0;
20'b00000010010000000010 : ColourData = 12'hDF0;
20'b00000010100000000010 : ColourData = 12'hDF0;
20'b00000010110000000010 : ColourData = 12'hDF0;
20'b00000011000000000010 : ColourData = 12'hDF0;
20'b00000011010000000010 : ColourData = 12'hDF0;
20'b00000011100000000010 : ColourData = 12'hDF0;
20'b00000011110000000010 : ColourData = 12'hDF0;
20'b00000100000000000010 : ColourData = 12'hDF0;
20'b00000100010000000010 : ColourData = 12'hDF0;
20'b00000100100000000010 : ColourData = 12'hFFF;
20'b00000100110000000010 : ColourData = 12'hFFF;
20'b00000101000000000010 : ColourData = 12'hFFF;
20'b00000101010000000010 : ColourData = 12'hFFF;
20'b00000101100000000010 : ColourData = 12'hFFF;
20'b00000101110000000010 : ColourData = 12'hFFF;
20'b00000110000000000010 : ColourData = 12'hFFF;
20'b00000000000000000011 : ColourData = 12'hFFF;
20'b00000000010000000011 : ColourData = 12'hFFF;
20'b00000000100000000011 : ColourData = 12'hFFF;
20'b00000000110000000011 : ColourData = 12'hFFF;
20'b00000001000000000011 : ColourData = 12'hFFF;
20'b00000001010000000011 : ColourData = 12'hFFF;
20'b00000001100000000011 : ColourData = 12'hDF0;
20'b00000001110000000011 : ColourData = 12'hDF0;
20'b00000010000000000011 : ColourData = 12'hDF0;
20'b00000010010000000011 : ColourData = 12'hDF0;
20'b00000010100000000011 : ColourData = 12'hDF0;
20'b00000010110000000011 : ColourData = 12'hDF0;
20'b00000011000000000011 : ColourData = 12'hDF0;
20'b00000011010000000011 : ColourData = 12'hDF0;
20'b00000011100000000011 : ColourData = 12'hDF0;
20'b00000011110000000011 : ColourData = 12'hDF0;
20'b00000100000000000011 : ColourData = 12'hDF0;
20'b00000100010000000011 : ColourData = 12'hDF0;
20'b00000100100000000011 : ColourData = 12'hDF0;
20'b00000100110000000011 : ColourData = 12'hFFF;
20'b00000101000000000011 : ColourData = 12'hFFF;
20'b00000101010000000011 : ColourData = 12'hFFF;
20'b00000101100000000011 : ColourData = 12'hFFF;
20'b00000101110000000011 : ColourData = 12'hFFF;
20'b00000110000000000011 : ColourData = 12'hFFF;
20'b00000000000000000100 : ColourData = 12'hFFF;
20'b00000000010000000100 : ColourData = 12'hFFF;
20'b00000000100000000100 : ColourData = 12'hFFF;
20'b00000000110000000100 : ColourData = 12'hFFF;
20'b00000001000000000100 : ColourData = 12'hDF0;
20'b00000001010000000100 : ColourData = 12'hDF0;
20'b00000001100000000100 : ColourData = 12'hDF0;
20'b00000001110000000100 : ColourData = 12'hDF0;
20'b00000010000000000100 : ColourData = 12'hDF0;
20'b00000010010000000100 : ColourData = 12'hDF0;
20'b00000010100000000100 : ColourData = 12'hDF0;
20'b00000010110000000100 : ColourData = 12'hDF0;
20'b00000011000000000100 : ColourData = 12'hDF0;
20'b00000011010000000100 : ColourData = 12'hDF0;
20'b00000011100000000100 : ColourData = 12'hDF0;
20'b00000011110000000100 : ColourData = 12'hDF0;
20'b00000100000000000100 : ColourData = 12'hDF0;
20'b00000100010000000100 : ColourData = 12'hDF0;
20'b00000100100000000100 : ColourData = 12'hDF0;
20'b00000100110000000100 : ColourData = 12'hDF0;
20'b00000101000000000100 : ColourData = 12'hDF0;
20'b00000101010000000100 : ColourData = 12'hFFF;
20'b00000101100000000100 : ColourData = 12'hFFF;
20'b00000101110000000100 : ColourData = 12'hFFF;
20'b00000110000000000100 : ColourData = 12'hFFF;
20'b00000000000000000101 : ColourData = 12'hFFF;
20'b00000000010000000101 : ColourData = 12'hFFF;
20'b00000000100000000101 : ColourData = 12'hFFF;
20'b00000000110000000101 : ColourData = 12'hFFF;
20'b00000001000000000101 : ColourData = 12'hDF0;
20'b00000001010000000101 : ColourData = 12'hDF0;
20'b00000001100000000101 : ColourData = 12'hDF0;
20'b00000001110000000101 : ColourData = 12'hDF0;
20'b00000010000000000101 : ColourData = 12'hDF0;
20'b00000010010000000101 : ColourData = 12'hDF0;
20'b00000010100000000101 : ColourData = 12'hDF0;
20'b00000010110000000101 : ColourData = 12'hDF0;
20'b00000011000000000101 : ColourData = 12'hDF0;
20'b00000011010000000101 : ColourData = 12'hDF0;
20'b00000011100000000101 : ColourData = 12'hDF0;
20'b00000011110000000101 : ColourData = 12'hDF0;
20'b00000100000000000101 : ColourData = 12'hDF0;
20'b00000100010000000101 : ColourData = 12'hDF0;
20'b00000100100000000101 : ColourData = 12'hDF0;
20'b00000100110000000101 : ColourData = 12'hDF0;
20'b00000101000000000101 : ColourData = 12'hDF0;
20'b00000101010000000101 : ColourData = 12'hFFF;
20'b00000101100000000101 : ColourData = 12'hFFF;
20'b00000101110000000101 : ColourData = 12'hFFF;
20'b00000110000000000101 : ColourData = 12'hFFF;
20'b00000000000000000110 : ColourData = 12'hFFF;
20'b00000000010000000110 : ColourData = 12'hFFF;
20'b00000000100000000110 : ColourData = 12'hFFF;
20'b00000000110000000110 : ColourData = 12'hDF0;
20'b00000001000000000110 : ColourData = 12'hDF0;
20'b00000001010000000110 : ColourData = 12'hDF0;
20'b00000001100000000110 : ColourData = 12'hDF0;
20'b00000001110000000110 : ColourData = 12'hDF0;
20'b00000010000000000110 : ColourData = 12'h000;
20'b00000010010000000110 : ColourData = 12'h000;
20'b00000010100000000110 : ColourData = 12'h000;
20'b00000010110000000110 : ColourData = 12'hDF0;
20'b00000011000000000110 : ColourData = 12'hDF0;
20'b00000011010000000110 : ColourData = 12'hDF0;
20'b00000011100000000110 : ColourData = 12'hDF0;
20'b00000011110000000110 : ColourData = 12'hDF0;
20'b00000100000000000110 : ColourData = 12'hDF0;
20'b00000100010000000110 : ColourData = 12'hDF0;
20'b00000100100000000110 : ColourData = 12'hDF0;
20'b00000100110000000110 : ColourData = 12'hDF0;
20'b00000101000000000110 : ColourData = 12'hFFF;
20'b00000101010000000110 : ColourData = 12'hFFF;
20'b00000101100000000110 : ColourData = 12'hFFF;
20'b00000101110000000110 : ColourData = 12'hFFF;
20'b00000110000000000110 : ColourData = 12'hFFF;
20'b00000000000000000111 : ColourData = 12'hFFF;
20'b00000000010000000111 : ColourData = 12'hFFF;
20'b00000000100000000111 : ColourData = 12'hDF0;
20'b00000000110000000111 : ColourData = 12'hDF0;
20'b00000001000000000111 : ColourData = 12'hDF0;
20'b00000001010000000111 : ColourData = 12'hDF0;
20'b00000001100000000111 : ColourData = 12'hDF0;
20'b00000001110000000111 : ColourData = 12'hDF0;
20'b00000010000000000111 : ColourData = 12'h000;
20'b00000010010000000111 : ColourData = 12'h000;
20'b00000010100000000111 : ColourData = 12'h000;
20'b00000010110000000111 : ColourData = 12'hDF0;
20'b00000011000000000111 : ColourData = 12'hDF0;
20'b00000011010000000111 : ColourData = 12'hDF0;
20'b00000011100000000111 : ColourData = 12'hDF0;
20'b00000011110000000111 : ColourData = 12'hDF0;
20'b00000100000000000111 : ColourData = 12'hDF0;
20'b00000100010000000111 : ColourData = 12'hDF0;
20'b00000100100000000111 : ColourData = 12'hDF0;
20'b00000100110000000111 : ColourData = 12'hFFF;
20'b00000101000000000111 : ColourData = 12'hFFF;
20'b00000101010000000111 : ColourData = 12'hFFF;
20'b00000101100000000111 : ColourData = 12'hFFF;
20'b00000101110000000111 : ColourData = 12'hFFF;
20'b00000110000000000111 : ColourData = 12'hFFF;
20'b00000000000000001000 : ColourData = 12'hFFF;
20'b00000000010000001000 : ColourData = 12'hFFF;
20'b00000000100000001000 : ColourData = 12'hDF0;
20'b00000000110000001000 : ColourData = 12'hDF0;
20'b00000001000000001000 : ColourData = 12'hDF0;
20'b00000001010000001000 : ColourData = 12'hDF0;
20'b00000001100000001000 : ColourData = 12'hDF0;
20'b00000001110000001000 : ColourData = 12'hDF0;
20'b00000010000000001000 : ColourData = 12'h000;
20'b00000010010000001000 : ColourData = 12'h000;
20'b00000010100000001000 : ColourData = 12'h000;
20'b00000010110000001000 : ColourData = 12'hDF0;
20'b00000011000000001000 : ColourData = 12'hDF0;
20'b00000011010000001000 : ColourData = 12'hDF0;
20'b00000011100000001000 : ColourData = 12'hDF0;
20'b00000011110000001000 : ColourData = 12'hDF0;
20'b00000100000000001000 : ColourData = 12'hDF0;
20'b00000100010000001000 : ColourData = 12'hDF0;
20'b00000100100000001000 : ColourData = 12'hFFF;
20'b00000100110000001000 : ColourData = 12'hFFF;
20'b00000101000000001000 : ColourData = 12'hFFF;
20'b00000101010000001000 : ColourData = 12'hFFF;
20'b00000101100000001000 : ColourData = 12'hFFF;
20'b00000101110000001000 : ColourData = 12'hFFF;
20'b00000110000000001000 : ColourData = 12'hFFF;
20'b00000000000000001001 : ColourData = 12'hFFF;
20'b00000000010000001001 : ColourData = 12'hDF0;
20'b00000000100000001001 : ColourData = 12'hDF0;
20'b00000000110000001001 : ColourData = 12'hDF0;
20'b00000001000000001001 : ColourData = 12'hDF0;
20'b00000001010000001001 : ColourData = 12'hDF0;
20'b00000001100000001001 : ColourData = 12'hDF0;
20'b00000001110000001001 : ColourData = 12'hDF0;
20'b00000010000000001001 : ColourData = 12'hDF0;
20'b00000010010000001001 : ColourData = 12'hDF0;
20'b00000010100000001001 : ColourData = 12'hDF0;
20'b00000010110000001001 : ColourData = 12'hDF0;
20'b00000011000000001001 : ColourData = 12'hDF0;
20'b00000011010000001001 : ColourData = 12'hDF0;
20'b00000011100000001001 : ColourData = 12'hDF0;
20'b00000011110000001001 : ColourData = 12'hDF0;
20'b00000100000000001001 : ColourData = 12'hDF0;
20'b00000100010000001001 : ColourData = 12'hFFF;
20'b00000100100000001001 : ColourData = 12'hFFF;
20'b00000100110000001001 : ColourData = 12'hFFF;
20'b00000101000000001001 : ColourData = 12'hFFF;
20'b00000101010000001001 : ColourData = 12'hFFF;
20'b00000101100000001001 : ColourData = 12'hFFF;
20'b00000101110000001001 : ColourData = 12'hFFF;
20'b00000110000000001001 : ColourData = 12'hFFF;
20'b00000000000000001010 : ColourData = 12'hFFF;
20'b00000000010000001010 : ColourData = 12'hDF0;
20'b00000000100000001010 : ColourData = 12'hDF0;
20'b00000000110000001010 : ColourData = 12'hDF0;
20'b00000001000000001010 : ColourData = 12'hDF0;
20'b00000001010000001010 : ColourData = 12'hDF0;
20'b00000001100000001010 : ColourData = 12'hDF0;
20'b00000001110000001010 : ColourData = 12'hDF0;
20'b00000010000000001010 : ColourData = 12'hDF0;
20'b00000010010000001010 : ColourData = 12'hDF0;
20'b00000010100000001010 : ColourData = 12'hDF0;
20'b00000010110000001010 : ColourData = 12'hDF0;
20'b00000011000000001010 : ColourData = 12'hDF0;
20'b00000011010000001010 : ColourData = 12'hDF0;
20'b00000011100000001010 : ColourData = 12'hDF0;
20'b00000011110000001010 : ColourData = 12'hDF0;
20'b00000100000000001010 : ColourData = 12'hFFF;
20'b00000100010000001010 : ColourData = 12'hFFF;
20'b00000100100000001010 : ColourData = 12'hFFF;
20'b00000100110000001010 : ColourData = 12'hFFF;
20'b00000101000000001010 : ColourData = 12'hFFF;
20'b00000101010000001010 : ColourData = 12'hFFF;
20'b00000101100000001010 : ColourData = 12'hFFF;
20'b00000101110000001010 : ColourData = 12'hFFF;
20'b00000110000000001010 : ColourData = 12'hFFF;
20'b00000000000000001011 : ColourData = 12'hFFF;
20'b00000000010000001011 : ColourData = 12'hDF0;
20'b00000000100000001011 : ColourData = 12'hDF0;
20'b00000000110000001011 : ColourData = 12'hDF0;
20'b00000001000000001011 : ColourData = 12'hDF0;
20'b00000001010000001011 : ColourData = 12'hDF0;
20'b00000001100000001011 : ColourData = 12'hDF0;
20'b00000001110000001011 : ColourData = 12'hDF0;
20'b00000010000000001011 : ColourData = 12'hDF0;
20'b00000010010000001011 : ColourData = 12'hDF0;
20'b00000010100000001011 : ColourData = 12'hDF0;
20'b00000010110000001011 : ColourData = 12'hDF0;
20'b00000011000000001011 : ColourData = 12'hDF0;
20'b00000011010000001011 : ColourData = 12'hDF0;
20'b00000011100000001011 : ColourData = 12'hDF0;
20'b00000011110000001011 : ColourData = 12'hFFF;
20'b00000100000000001011 : ColourData = 12'hFFF;
20'b00000100010000001011 : ColourData = 12'hFFF;
20'b00000100100000001011 : ColourData = 12'hFFF;
20'b00000100110000001011 : ColourData = 12'hFFF;
20'b00000101000000001011 : ColourData = 12'hFFF;
20'b00000101010000001011 : ColourData = 12'hFFF;
20'b00000101100000001011 : ColourData = 12'hFFF;
20'b00000101110000001011 : ColourData = 12'hFFF;
20'b00000110000000001011 : ColourData = 12'hFFF;
20'b00000000000000001100 : ColourData = 12'hFFF;
20'b00000000010000001100 : ColourData = 12'hDF0;
20'b00000000100000001100 : ColourData = 12'hDF0;
20'b00000000110000001100 : ColourData = 12'hDF0;
20'b00000001000000001100 : ColourData = 12'hDF0;
20'b00000001010000001100 : ColourData = 12'hDF0;
20'b00000001100000001100 : ColourData = 12'hDF0;
20'b00000001110000001100 : ColourData = 12'hDF0;
20'b00000010000000001100 : ColourData = 12'hDF0;
20'b00000010010000001100 : ColourData = 12'hDF0;
20'b00000010100000001100 : ColourData = 12'hDF0;
20'b00000010110000001100 : ColourData = 12'hDF0;
20'b00000011000000001100 : ColourData = 12'hDF0;
20'b00000011010000001100 : ColourData = 12'hDF0;
20'b00000011100000001100 : ColourData = 12'hFFF;
20'b00000011110000001100 : ColourData = 12'hFFF;
20'b00000100000000001100 : ColourData = 12'hFFF;
20'b00000100010000001100 : ColourData = 12'hFFF;
20'b00000100100000001100 : ColourData = 12'hFFF;
20'b00000100110000001100 : ColourData = 12'hFFF;
20'b00000101000000001100 : ColourData = 12'hFFF;
20'b00000101010000001100 : ColourData = 12'hFFF;
20'b00000101100000001100 : ColourData = 12'hFFF;
20'b00000101110000001100 : ColourData = 12'hFFF;
20'b00000110000000001100 : ColourData = 12'hFFF;
20'b00000000000000001101 : ColourData = 12'hFFF;
20'b00000000010000001101 : ColourData = 12'hDF0;
20'b00000000100000001101 : ColourData = 12'hDF0;
20'b00000000110000001101 : ColourData = 12'hDF0;
20'b00000001000000001101 : ColourData = 12'hDF0;
20'b00000001010000001101 : ColourData = 12'hDF0;
20'b00000001100000001101 : ColourData = 12'hDF0;
20'b00000001110000001101 : ColourData = 12'hDF0;
20'b00000010000000001101 : ColourData = 12'hDF0;
20'b00000010010000001101 : ColourData = 12'hDF0;
20'b00000010100000001101 : ColourData = 12'hDF0;
20'b00000010110000001101 : ColourData = 12'hDF0;
20'b00000011000000001101 : ColourData = 12'hDF0;
20'b00000011010000001101 : ColourData = 12'hDF0;
20'b00000011100000001101 : ColourData = 12'hDF0;
20'b00000011110000001101 : ColourData = 12'hFFF;
20'b00000100000000001101 : ColourData = 12'hFFF;
20'b00000100010000001101 : ColourData = 12'hFFF;
20'b00000100100000001101 : ColourData = 12'hFFF;
20'b00000100110000001101 : ColourData = 12'hFFF;
20'b00000101000000001101 : ColourData = 12'hFFF;
20'b00000101010000001101 : ColourData = 12'hFFF;
20'b00000101100000001101 : ColourData = 12'hFFF;
20'b00000101110000001101 : ColourData = 12'hFFF;
20'b00000110000000001101 : ColourData = 12'hFFF;
20'b00000000000000001110 : ColourData = 12'hFFF;
20'b00000000010000001110 : ColourData = 12'hDF0;
20'b00000000100000001110 : ColourData = 12'hDF0;
20'b00000000110000001110 : ColourData = 12'hDF0;
20'b00000001000000001110 : ColourData = 12'hDF0;
20'b00000001010000001110 : ColourData = 12'hDF0;
20'b00000001100000001110 : ColourData = 12'hDF0;
20'b00000001110000001110 : ColourData = 12'hDF0;
20'b00000010000000001110 : ColourData = 12'hDF0;
20'b00000010010000001110 : ColourData = 12'hDF0;
20'b00000010100000001110 : ColourData = 12'hDF0;
20'b00000010110000001110 : ColourData = 12'hDF0;
20'b00000011000000001110 : ColourData = 12'hDF0;
20'b00000011010000001110 : ColourData = 12'hDF0;
20'b00000011100000001110 : ColourData = 12'hDF0;
20'b00000011110000001110 : ColourData = 12'hDF0;
20'b00000100000000001110 : ColourData = 12'hFFF;
20'b00000100010000001110 : ColourData = 12'hFFF;
20'b00000100100000001110 : ColourData = 12'hFFF;
20'b00000100110000001110 : ColourData = 12'hFFF;
20'b00000101000000001110 : ColourData = 12'hFFF;
20'b00000101010000001110 : ColourData = 12'hFFF;
20'b00000101100000001110 : ColourData = 12'hFFF;
20'b00000101110000001110 : ColourData = 12'hFFF;
20'b00000110000000001110 : ColourData = 12'hFFF;
20'b00000000000000001111 : ColourData = 12'hFFF;
20'b00000000010000001111 : ColourData = 12'hDF0;
20'b00000000100000001111 : ColourData = 12'hDF0;
20'b00000000110000001111 : ColourData = 12'hDF0;
20'b00000001000000001111 : ColourData = 12'hDF0;
20'b00000001010000001111 : ColourData = 12'hDF0;
20'b00000001100000001111 : ColourData = 12'hDF0;
20'b00000001110000001111 : ColourData = 12'hDF0;
20'b00000010000000001111 : ColourData = 12'hDF0;
20'b00000010010000001111 : ColourData = 12'hDF0;
20'b00000010100000001111 : ColourData = 12'hDF0;
20'b00000010110000001111 : ColourData = 12'hDF0;
20'b00000011000000001111 : ColourData = 12'hDF0;
20'b00000011010000001111 : ColourData = 12'hDF0;
20'b00000011100000001111 : ColourData = 12'hDF0;
20'b00000011110000001111 : ColourData = 12'hDF0;
20'b00000100000000001111 : ColourData = 12'hDF0;
20'b00000100010000001111 : ColourData = 12'hFFF;
20'b00000100100000001111 : ColourData = 12'hFFF;
20'b00000100110000001111 : ColourData = 12'hFFF;
20'b00000101000000001111 : ColourData = 12'hFFF;
20'b00000101010000001111 : ColourData = 12'hFFF;
20'b00000101100000001111 : ColourData = 12'hFFF;
20'b00000101110000001111 : ColourData = 12'hFFF;
20'b00000110000000001111 : ColourData = 12'hFFF;
20'b00000000000000010000 : ColourData = 12'hFFF;
20'b00000000010000010000 : ColourData = 12'hFFF;
20'b00000000100000010000 : ColourData = 12'hDF0;
20'b00000000110000010000 : ColourData = 12'hDF0;
20'b00000001000000010000 : ColourData = 12'hDF0;
20'b00000001010000010000 : ColourData = 12'hDF0;
20'b00000001100000010000 : ColourData = 12'hDF0;
20'b00000001110000010000 : ColourData = 12'hDF0;
20'b00000010000000010000 : ColourData = 12'hDF0;
20'b00000010010000010000 : ColourData = 12'hDF0;
20'b00000010100000010000 : ColourData = 12'hDF0;
20'b00000010110000010000 : ColourData = 12'hDF0;
20'b00000011000000010000 : ColourData = 12'hDF0;
20'b00000011010000010000 : ColourData = 12'hDF0;
20'b00000011100000010000 : ColourData = 12'hDF0;
20'b00000011110000010000 : ColourData = 12'hDF0;
20'b00000100000000010000 : ColourData = 12'hDF0;
20'b00000100010000010000 : ColourData = 12'hDF0;
20'b00000100100000010000 : ColourData = 12'hFFF;
20'b00000100110000010000 : ColourData = 12'hFFF;
20'b00000101000000010000 : ColourData = 12'hFFF;
20'b00000101010000010000 : ColourData = 12'hFFF;
20'b00000101100000010000 : ColourData = 12'hFFF;
20'b00000101110000010000 : ColourData = 12'hFFF;
20'b00000110000000010000 : ColourData = 12'hFFF;
20'b00000000000000010001 : ColourData = 12'hFFF;
20'b00000000010000010001 : ColourData = 12'hFFF;
20'b00000000100000010001 : ColourData = 12'hDF0;
20'b00000000110000010001 : ColourData = 12'hDF0;
20'b00000001000000010001 : ColourData = 12'hDF0;
20'b00000001010000010001 : ColourData = 12'hDF0;
20'b00000001100000010001 : ColourData = 12'hDF0;
20'b00000001110000010001 : ColourData = 12'hDF0;
20'b00000010000000010001 : ColourData = 12'hDF0;
20'b00000010010000010001 : ColourData = 12'hDF0;
20'b00000010100000010001 : ColourData = 12'hDF0;
20'b00000010110000010001 : ColourData = 12'hDF0;
20'b00000011000000010001 : ColourData = 12'hDF0;
20'b00000011010000010001 : ColourData = 12'hDF0;
20'b00000011100000010001 : ColourData = 12'hDF0;
20'b00000011110000010001 : ColourData = 12'hDF0;
20'b00000100000000010001 : ColourData = 12'hDF0;
20'b00000100010000010001 : ColourData = 12'hDF0;
20'b00000100100000010001 : ColourData = 12'hDF0;
20'b00000100110000010001 : ColourData = 12'hFFF;
20'b00000101000000010001 : ColourData = 12'hFFF;
20'b00000101010000010001 : ColourData = 12'hFFF;
20'b00000101100000010001 : ColourData = 12'hFFF;
20'b00000101110000010001 : ColourData = 12'hFFF;
20'b00000110000000010001 : ColourData = 12'hFFF;
20'b00000000000000010010 : ColourData = 12'hFFF;
20'b00000000010000010010 : ColourData = 12'hFFF;
20'b00000000100000010010 : ColourData = 12'hFFF;
20'b00000000110000010010 : ColourData = 12'hDF0;
20'b00000001000000010010 : ColourData = 12'hDF0;
20'b00000001010000010010 : ColourData = 12'hDF0;
20'b00000001100000010010 : ColourData = 12'hDF0;
20'b00000001110000010010 : ColourData = 12'hDF0;
20'b00000010000000010010 : ColourData = 12'hDF0;
20'b00000010010000010010 : ColourData = 12'hDF0;
20'b00000010100000010010 : ColourData = 12'hDF0;
20'b00000010110000010010 : ColourData = 12'hDF0;
20'b00000011000000010010 : ColourData = 12'hDF0;
20'b00000011010000010010 : ColourData = 12'hDF0;
20'b00000011100000010010 : ColourData = 12'hDF0;
20'b00000011110000010010 : ColourData = 12'hDF0;
20'b00000100000000010010 : ColourData = 12'hDF0;
20'b00000100010000010010 : ColourData = 12'hDF0;
20'b00000100100000010010 : ColourData = 12'hDF0;
20'b00000100110000010010 : ColourData = 12'hDF0;
20'b00000101000000010010 : ColourData = 12'hFFF;
20'b00000101010000010010 : ColourData = 12'hFFF;
20'b00000101100000010010 : ColourData = 12'hFFF;
20'b00000101110000010010 : ColourData = 12'hFFF;
20'b00000110000000010010 : ColourData = 12'hFFF;
20'b00000000000000010011 : ColourData = 12'hFFF;
20'b00000000010000010011 : ColourData = 12'hFFF;
20'b00000000100000010011 : ColourData = 12'hFFF;
20'b00000000110000010011 : ColourData = 12'hFFF;
20'b00000001000000010011 : ColourData = 12'hDF0;
20'b00000001010000010011 : ColourData = 12'hDF0;
20'b00000001100000010011 : ColourData = 12'hDF0;
20'b00000001110000010011 : ColourData = 12'hDF0;
20'b00000010000000010011 : ColourData = 12'hDF0;
20'b00000010010000010011 : ColourData = 12'hDF0;
20'b00000010100000010011 : ColourData = 12'hDF0;
20'b00000010110000010011 : ColourData = 12'hDF0;
20'b00000011000000010011 : ColourData = 12'hDF0;
20'b00000011010000010011 : ColourData = 12'hDF0;
20'b00000011100000010011 : ColourData = 12'hDF0;
20'b00000011110000010011 : ColourData = 12'hDF0;
20'b00000100000000010011 : ColourData = 12'hDF0;
20'b00000100010000010011 : ColourData = 12'hDF0;
20'b00000100100000010011 : ColourData = 12'hDF0;
20'b00000100110000010011 : ColourData = 12'hDF0;
20'b00000101000000010011 : ColourData = 12'hDF0;
20'b00000101010000010011 : ColourData = 12'hFFF;
20'b00000101100000010011 : ColourData = 12'hFFF;
20'b00000101110000010011 : ColourData = 12'hFFF;
20'b00000110000000010011 : ColourData = 12'hFFF;
20'b00000000000000010100 : ColourData = 12'hFFF;
20'b00000000010000010100 : ColourData = 12'hFFF;
20'b00000000100000010100 : ColourData = 12'hFFF;
20'b00000000110000010100 : ColourData = 12'hFFF;
20'b00000001000000010100 : ColourData = 12'hDF0;
20'b00000001010000010100 : ColourData = 12'hDF0;
20'b00000001100000010100 : ColourData = 12'hDF0;
20'b00000001110000010100 : ColourData = 12'hDF0;
20'b00000010000000010100 : ColourData = 12'hDF0;
20'b00000010010000010100 : ColourData = 12'hDF0;
20'b00000010100000010100 : ColourData = 12'hDF0;
20'b00000010110000010100 : ColourData = 12'hDF0;
20'b00000011000000010100 : ColourData = 12'hDF0;
20'b00000011010000010100 : ColourData = 12'hDF0;
20'b00000011100000010100 : ColourData = 12'hDF0;
20'b00000011110000010100 : ColourData = 12'hDF0;
20'b00000100000000010100 : ColourData = 12'hDF0;
20'b00000100010000010100 : ColourData = 12'hDF0;
20'b00000100100000010100 : ColourData = 12'hDF0;
20'b00000100110000010100 : ColourData = 12'hDF0;
20'b00000101000000010100 : ColourData = 12'hDF0;
20'b00000101010000010100 : ColourData = 12'hFFF;
20'b00000101100000010100 : ColourData = 12'hFFF;
20'b00000101110000010100 : ColourData = 12'hFFF;
20'b00000110000000010100 : ColourData = 12'hFFF;
20'b00000000000000010101 : ColourData = 12'hFFF;
20'b00000000010000010101 : ColourData = 12'hFFF;
20'b00000000100000010101 : ColourData = 12'hFFF;
20'b00000000110000010101 : ColourData = 12'hFFF;
20'b00000001000000010101 : ColourData = 12'hFFF;
20'b00000001010000010101 : ColourData = 12'hFFF;
20'b00000001100000010101 : ColourData = 12'hDF0;
20'b00000001110000010101 : ColourData = 12'hDF0;
20'b00000010000000010101 : ColourData = 12'hDF0;
20'b00000010010000010101 : ColourData = 12'hDF0;
20'b00000010100000010101 : ColourData = 12'hDF0;
20'b00000010110000010101 : ColourData = 12'hDF0;
20'b00000011000000010101 : ColourData = 12'hDF0;
20'b00000011010000010101 : ColourData = 12'hDF0;
20'b00000011100000010101 : ColourData = 12'hDF0;
20'b00000011110000010101 : ColourData = 12'hDF0;
20'b00000100000000010101 : ColourData = 12'hDF0;
20'b00000100010000010101 : ColourData = 12'hDF0;
20'b00000100100000010101 : ColourData = 12'hDF0;
20'b00000100110000010101 : ColourData = 12'hFFF;
20'b00000101000000010101 : ColourData = 12'hFFF;
20'b00000101010000010101 : ColourData = 12'hFFF;
20'b00000101100000010101 : ColourData = 12'hFFF;
20'b00000101110000010101 : ColourData = 12'hFFF;
20'b00000110000000010101 : ColourData = 12'hFFF;
20'b00000000000000010110 : ColourData = 12'hFFF;
20'b00000000010000010110 : ColourData = 12'hFFF;
20'b00000000100000010110 : ColourData = 12'hFFF;
20'b00000000110000010110 : ColourData = 12'hFFF;
20'b00000001000000010110 : ColourData = 12'hFFF;
20'b00000001010000010110 : ColourData = 12'hFFF;
20'b00000001100000010110 : ColourData = 12'hFFF;
20'b00000001110000010110 : ColourData = 12'hDF0;
20'b00000010000000010110 : ColourData = 12'hDF0;
20'b00000010010000010110 : ColourData = 12'hDF0;
20'b00000010100000010110 : ColourData = 12'hDF0;
20'b00000010110000010110 : ColourData = 12'hDF0;
20'b00000011000000010110 : ColourData = 12'hDF0;
20'b00000011010000010110 : ColourData = 12'hDF0;
20'b00000011100000010110 : ColourData = 12'hDF0;
20'b00000011110000010110 : ColourData = 12'hDF0;
20'b00000100000000010110 : ColourData = 12'hDF0;
20'b00000100010000010110 : ColourData = 12'hDF0;
20'b00000100100000010110 : ColourData = 12'hFFF;
20'b00000100110000010110 : ColourData = 12'hFFF;
20'b00000101000000010110 : ColourData = 12'hFFF;
20'b00000101010000010110 : ColourData = 12'hFFF;
20'b00000101100000010110 : ColourData = 12'hFFF;
20'b00000101110000010110 : ColourData = 12'hFFF;
20'b00000110000000010110 : ColourData = 12'hFFF;
20'b00000000000000010111 : ColourData = 12'hFFF;
20'b00000000010000010111 : ColourData = 12'hFFF;
20'b00000000100000010111 : ColourData = 12'hFFF;
20'b00000000110000010111 : ColourData = 12'hFFF;
20'b00000001000000010111 : ColourData = 12'hFFF;
20'b00000001010000010111 : ColourData = 12'hFFF;
20'b00000001100000010111 : ColourData = 12'hFFF;
20'b00000001110000010111 : ColourData = 12'hFFF;
20'b00000010000000010111 : ColourData = 12'hFFF;
20'b00000010010000010111 : ColourData = 12'hDF0;
20'b00000010100000010111 : ColourData = 12'hDF0;
20'b00000010110000010111 : ColourData = 12'hDF0;
20'b00000011000000010111 : ColourData = 12'hDF0;
20'b00000011010000010111 : ColourData = 12'hDF0;
20'b00000011100000010111 : ColourData = 12'hDF0;
20'b00000011110000010111 : ColourData = 12'hDF0;
20'b00000100000000010111 : ColourData = 12'hFFF;
20'b00000100010000010111 : ColourData = 12'hFFF;
20'b00000100100000010111 : ColourData = 12'hFFF;
20'b00000100110000010111 : ColourData = 12'hFFF;
20'b00000101000000010111 : ColourData = 12'hFFF;
20'b00000101010000010111 : ColourData = 12'hFFF;
20'b00000101100000010111 : ColourData = 12'hFFF;
20'b00000101110000010111 : ColourData = 12'hFFF;
20'b00000110000000010111 : ColourData = 12'hFFF;
20'b00000000000000011000 : ColourData = 12'hFFF;
20'b00000000010000011000 : ColourData = 12'hFFF;
20'b00000000100000011000 : ColourData = 12'hFFF;
20'b00000000110000011000 : ColourData = 12'hFFF;
20'b00000001000000011000 : ColourData = 12'hFFF;
20'b00000001010000011000 : ColourData = 12'hFFF;
20'b00000001100000011000 : ColourData = 12'hFFF;
20'b00000001110000011000 : ColourData = 12'hFFF;
20'b00000010000000011000 : ColourData = 12'hFFF;
20'b00000010010000011000 : ColourData = 12'hFFF;
20'b00000010100000011000 : ColourData = 12'hFFF;
20'b00000010110000011000 : ColourData = 12'hFFF;
20'b00000011000000011000 : ColourData = 12'hFFF;
20'b00000011010000011000 : ColourData = 12'hFFF;
20'b00000011100000011000 : ColourData = 12'hFFF;
20'b00000011110000011000 : ColourData = 12'hFFF;
20'b00000100000000011000 : ColourData = 12'hFFF;
20'b00000100010000011000 : ColourData = 12'hFFF;
20'b00000100100000011000 : ColourData = 12'hFFF;
20'b00000100110000011000 : ColourData = 12'hFFF;
20'b00000101000000011000 : ColourData = 12'hFFF;
20'b00000101010000011000 : ColourData = 12'hFFF;
20'b00000101100000011000 : ColourData = 12'hFFF;
20'b00000101110000011000 : ColourData = 12'hFFF;
20'b00000110000000011000 : ColourData = 12'hFFF;

    
default: ColourData = 12'h000;

endcase
end

endmodule