module TankImage(

  input Master_Clock_In,
  input [9 : 0] xInput,
  input [9 : 0] yInput,
  output reg [11:0] ColourData = 12'h000

);

(* rom_style = "block" *)

reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

always @(posedge Master_Clock_In)
begin
  a = xInput % 60;
  b = yInput % 60;

Inputs = {a, b};

    case(Inputs)
    
    
20'b00000000000000000000 : ColourData = 12'hFFF;
20'b00000000010000000000 : ColourData = 12'hFFF;
20'b00000000100000000000 : ColourData = 12'hFFF;
20'b00000000110000000000 : ColourData = 12'hFFF;
20'b00000001000000000000 : ColourData = 12'hFFF;
20'b00000001010000000000 : ColourData = 12'hFFF;
20'b00000001100000000000 : ColourData = 12'hFFF;
20'b00000001110000000000 : ColourData = 12'hFFF;
20'b00000010000000000000 : ColourData = 12'hFFF;
20'b00000010010000000000 : ColourData = 12'hFFF;
20'b00000010100000000000 : ColourData = 12'hFFF;
20'b00000010110000000000 : ColourData = 12'hFFF;
20'b00000011000000000000 : ColourData = 12'hFFF;
20'b00000011010000000000 : ColourData = 12'hFFF;
20'b00000011100000000000 : ColourData = 12'hFFF;
20'b00000011110000000000 : ColourData = 12'hFFF;
20'b00000100000000000000 : ColourData = 12'hFFF;
20'b00000100010000000000 : ColourData = 12'hFFF;
20'b00000100100000000000 : ColourData = 12'hFFF;
20'b00000100110000000000 : ColourData = 12'hFFF;
20'b00000101000000000000 : ColourData = 12'hFFF;
20'b00000101010000000000 : ColourData = 12'hFFF;
20'b00000101100000000000 : ColourData = 12'hFFF;
20'b00000101110000000000 : ColourData = 12'hFFF;
20'b00000110000000000000 : ColourData = 12'hFFF;
20'b00000110010000000000 : ColourData = 12'hFFF;
20'b00000110100000000000 : ColourData = 12'hFFF;
20'b00000110110000000000 : ColourData = 12'hAAA;
20'b00000111000000000000 : ColourData = 12'h000;
20'b00000111010000000000 : ColourData = 12'h000;
20'b00000111100000000000 : ColourData = 12'h000;
20'b00000111110000000000 : ColourData = 12'h000;
20'b00001000000000000000 : ColourData = 12'hAAA;
20'b00001000010000000000 : ColourData = 12'hFFF;
20'b00001000100000000000 : ColourData = 12'hFFF;
20'b00001000110000000000 : ColourData = 12'hFFF;
20'b00001001000000000000 : ColourData = 12'hFFF;
20'b00001001010000000000 : ColourData = 12'hFFF;
20'b00001001100000000000 : ColourData = 12'hFFF;
20'b00001001110000000000 : ColourData = 12'hFFF;
20'b00001010000000000000 : ColourData = 12'hFFF;
20'b00001010010000000000 : ColourData = 12'hFFF;
20'b00001010100000000000 : ColourData = 12'hFFF;
20'b00001010110000000000 : ColourData = 12'hFFF;
20'b00001011000000000000 : ColourData = 12'hFFF;
20'b00001011010000000000 : ColourData = 12'hFFF;
20'b00001011100000000000 : ColourData = 12'hFFF;
20'b00001011110000000000 : ColourData = 12'hFFF;
20'b00001100000000000000 : ColourData = 12'hFFF;
20'b00001100010000000000 : ColourData = 12'hFFF;
20'b00001100100000000000 : ColourData = 12'hFFF;
20'b00001100110000000000 : ColourData = 12'hFFF;
20'b00001101000000000000 : ColourData = 12'hFFF;
20'b00001101010000000000 : ColourData = 12'hFFF;
20'b00001101100000000000 : ColourData = 12'hFFF;
20'b00001101110000000000 : ColourData = 12'hFFF;
20'b00001110000000000000 : ColourData = 12'hFFF;
20'b00001110010000000000 : ColourData = 12'hFFF;
20'b00001110100000000000 : ColourData = 12'hFFF;
20'b00001110110000000000 : ColourData = 12'hFFF;
20'b00000000000000000001 : ColourData = 12'hFFF;
20'b00000000010000000001 : ColourData = 12'hFFF;
20'b00000000100000000001 : ColourData = 12'hFFF;
20'b00000000110000000001 : ColourData = 12'hFFF;
20'b00000001000000000001 : ColourData = 12'hFFF;
20'b00000001010000000001 : ColourData = 12'hFFF;
20'b00000001100000000001 : ColourData = 12'hFFF;
20'b00000001110000000001 : ColourData = 12'hFFF;
20'b00000010000000000001 : ColourData = 12'hFFF;
20'b00000010010000000001 : ColourData = 12'hFFF;
20'b00000010100000000001 : ColourData = 12'hFFF;
20'b00000010110000000001 : ColourData = 12'hFFF;
20'b00000011000000000001 : ColourData = 12'hFFF;
20'b00000011010000000001 : ColourData = 12'hFFF;
20'b00000011100000000001 : ColourData = 12'hFFF;
20'b00000011110000000001 : ColourData = 12'hFFF;
20'b00000100000000000001 : ColourData = 12'hFFF;
20'b00000100010000000001 : ColourData = 12'hFFF;
20'b00000100100000000001 : ColourData = 12'hFFF;
20'b00000100110000000001 : ColourData = 12'hFFF;
20'b00000101000000000001 : ColourData = 12'hFFF;
20'b00000101010000000001 : ColourData = 12'hFFF;
20'b00000101100000000001 : ColourData = 12'hFFF;
20'b00000101110000000001 : ColourData = 12'hFFF;
20'b00000110000000000001 : ColourData = 12'hFFF;
20'b00000110010000000001 : ColourData = 12'hFFF;
20'b00000110100000000001 : ColourData = 12'hFFF;
20'b00000110110000000001 : ColourData = 12'hAAA;
20'b00000111000000000001 : ColourData = 12'h000;
20'b00000111010000000001 : ColourData = 12'h000;
20'b00000111100000000001 : ColourData = 12'h000;
20'b00000111110000000001 : ColourData = 12'h000;
20'b00001000000000000001 : ColourData = 12'hAAA;
20'b00001000010000000001 : ColourData = 12'hFFF;
20'b00001000100000000001 : ColourData = 12'hFFF;
20'b00001000110000000001 : ColourData = 12'hFFF;
20'b00001001000000000001 : ColourData = 12'hFFF;
20'b00001001010000000001 : ColourData = 12'hFFF;
20'b00001001100000000001 : ColourData = 12'hFFF;
20'b00001001110000000001 : ColourData = 12'hFFF;
20'b00001010000000000001 : ColourData = 12'hFFF;
20'b00001010010000000001 : ColourData = 12'hFFF;
20'b00001010100000000001 : ColourData = 12'hFFF;
20'b00001010110000000001 : ColourData = 12'hFFF;
20'b00001011000000000001 : ColourData = 12'hFFF;
20'b00001011010000000001 : ColourData = 12'hFFF;
20'b00001011100000000001 : ColourData = 12'hFFF;
20'b00001011110000000001 : ColourData = 12'hFFF;
20'b00001100000000000001 : ColourData = 12'hFFF;
20'b00001100010000000001 : ColourData = 12'hFFF;
20'b00001100100000000001 : ColourData = 12'hFFF;
20'b00001100110000000001 : ColourData = 12'hFFF;
20'b00001101000000000001 : ColourData = 12'hFFF;
20'b00001101010000000001 : ColourData = 12'hFFF;
20'b00001101100000000001 : ColourData = 12'hFFF;
20'b00001101110000000001 : ColourData = 12'hFFF;
20'b00001110000000000001 : ColourData = 12'hFFF;
20'b00001110010000000001 : ColourData = 12'hFFF;
20'b00001110100000000001 : ColourData = 12'hFFF;
20'b00001110110000000001 : ColourData = 12'hFFF;
20'b00000000000000000010 : ColourData = 12'hFFF;
20'b00000000010000000010 : ColourData = 12'hFFF;
20'b00000000100000000010 : ColourData = 12'hFFF;
20'b00000000110000000010 : ColourData = 12'hFFF;
20'b00000001000000000010 : ColourData = 12'hFFF;
20'b00000001010000000010 : ColourData = 12'hFFF;
20'b00000001100000000010 : ColourData = 12'hFFF;
20'b00000001110000000010 : ColourData = 12'hFFF;
20'b00000010000000000010 : ColourData = 12'hFFF;
20'b00000010010000000010 : ColourData = 12'hFFF;
20'b00000010100000000010 : ColourData = 12'hFFF;
20'b00000010110000000010 : ColourData = 12'hFFF;
20'b00000011000000000010 : ColourData = 12'hFFF;
20'b00000011010000000010 : ColourData = 12'hFFF;
20'b00000011100000000010 : ColourData = 12'hFFF;
20'b00000011110000000010 : ColourData = 12'hFFF;
20'b00000100000000000010 : ColourData = 12'hFFF;
20'b00000100010000000010 : ColourData = 12'hFFF;
20'b00000100100000000010 : ColourData = 12'hFFF;
20'b00000100110000000010 : ColourData = 12'hFFF;
20'b00000101000000000010 : ColourData = 12'hFFF;
20'b00000101010000000010 : ColourData = 12'hFFF;
20'b00000101100000000010 : ColourData = 12'hFFF;
20'b00000101110000000010 : ColourData = 12'hFFF;
20'b00000110000000000010 : ColourData = 12'hFFF;
20'b00000110010000000010 : ColourData = 12'hFFF;
20'b00000110100000000010 : ColourData = 12'hFFF;
20'b00000110110000000010 : ColourData = 12'hAAA;
20'b00000111000000000010 : ColourData = 12'h000;
20'b00000111010000000010 : ColourData = 12'h000;
20'b00000111100000000010 : ColourData = 12'h000;
20'b00000111110000000010 : ColourData = 12'h000;
20'b00001000000000000010 : ColourData = 12'hAAA;
20'b00001000010000000010 : ColourData = 12'hFFF;
20'b00001000100000000010 : ColourData = 12'hFFF;
20'b00001000110000000010 : ColourData = 12'hFFF;
20'b00001001000000000010 : ColourData = 12'hFFF;
20'b00001001010000000010 : ColourData = 12'hFFF;
20'b00001001100000000010 : ColourData = 12'hFFF;
20'b00001001110000000010 : ColourData = 12'hFFF;
20'b00001010000000000010 : ColourData = 12'hFFF;
20'b00001010010000000010 : ColourData = 12'hFFF;
20'b00001010100000000010 : ColourData = 12'hFFF;
20'b00001010110000000010 : ColourData = 12'hFFF;
20'b00001011000000000010 : ColourData = 12'hFFF;
20'b00001011010000000010 : ColourData = 12'hFFF;
20'b00001011100000000010 : ColourData = 12'hFFF;
20'b00001011110000000010 : ColourData = 12'hFFF;
20'b00001100000000000010 : ColourData = 12'hFFF;
20'b00001100010000000010 : ColourData = 12'hFFF;
20'b00001100100000000010 : ColourData = 12'hFFF;
20'b00001100110000000010 : ColourData = 12'hFFF;
20'b00001101000000000010 : ColourData = 12'hFFF;
20'b00001101010000000010 : ColourData = 12'hFFF;
20'b00001101100000000010 : ColourData = 12'hFFF;
20'b00001101110000000010 : ColourData = 12'hFFF;
20'b00001110000000000010 : ColourData = 12'hFFF;
20'b00001110010000000010 : ColourData = 12'hFFF;
20'b00001110100000000010 : ColourData = 12'hFFF;
20'b00001110110000000010 : ColourData = 12'hFFF;
20'b00000000000000000011 : ColourData = 12'hFFF;
20'b00000000010000000011 : ColourData = 12'hFFF;
20'b00000000100000000011 : ColourData = 12'hFFF;
20'b00000000110000000011 : ColourData = 12'hFFF;
20'b00000001000000000011 : ColourData = 12'hFFF;
20'b00000001010000000011 : ColourData = 12'hFFF;
20'b00000001100000000011 : ColourData = 12'hFFF;
20'b00000001110000000011 : ColourData = 12'hFFF;
20'b00000010000000000011 : ColourData = 12'hFFF;
20'b00000010010000000011 : ColourData = 12'hFFF;
20'b00000010100000000011 : ColourData = 12'hFFF;
20'b00000010110000000011 : ColourData = 12'hFFF;
20'b00000011000000000011 : ColourData = 12'hFFF;
20'b00000011010000000011 : ColourData = 12'hFFF;
20'b00000011100000000011 : ColourData = 12'hFFF;
20'b00000011110000000011 : ColourData = 12'hFFF;
20'b00000100000000000011 : ColourData = 12'hFFF;
20'b00000100010000000011 : ColourData = 12'hFFF;
20'b00000100100000000011 : ColourData = 12'hFFF;
20'b00000100110000000011 : ColourData = 12'hFFF;
20'b00000101000000000011 : ColourData = 12'hFFF;
20'b00000101010000000011 : ColourData = 12'hFFF;
20'b00000101100000000011 : ColourData = 12'hFFF;
20'b00000101110000000011 : ColourData = 12'hFFF;
20'b00000110000000000011 : ColourData = 12'hFFF;
20'b00000110010000000011 : ColourData = 12'hFFF;
20'b00000110100000000011 : ColourData = 12'hFFF;
20'b00000110110000000011 : ColourData = 12'hAAA;
20'b00000111000000000011 : ColourData = 12'h000;
20'b00000111010000000011 : ColourData = 12'h000;
20'b00000111100000000011 : ColourData = 12'h000;
20'b00000111110000000011 : ColourData = 12'h000;
20'b00001000000000000011 : ColourData = 12'hAAA;
20'b00001000010000000011 : ColourData = 12'hFFF;
20'b00001000100000000011 : ColourData = 12'hFFF;
20'b00001000110000000011 : ColourData = 12'hFFF;
20'b00001001000000000011 : ColourData = 12'hFFF;
20'b00001001010000000011 : ColourData = 12'hFFF;
20'b00001001100000000011 : ColourData = 12'hFFF;
20'b00001001110000000011 : ColourData = 12'hFFF;
20'b00001010000000000011 : ColourData = 12'hFFF;
20'b00001010010000000011 : ColourData = 12'hFFF;
20'b00001010100000000011 : ColourData = 12'hFFF;
20'b00001010110000000011 : ColourData = 12'hFFF;
20'b00001011000000000011 : ColourData = 12'hFFF;
20'b00001011010000000011 : ColourData = 12'hFFF;
20'b00001011100000000011 : ColourData = 12'hFFF;
20'b00001011110000000011 : ColourData = 12'hFFF;
20'b00001100000000000011 : ColourData = 12'hFFF;
20'b00001100010000000011 : ColourData = 12'hFFF;
20'b00001100100000000011 : ColourData = 12'hFFF;
20'b00001100110000000011 : ColourData = 12'hFFF;
20'b00001101000000000011 : ColourData = 12'hFFF;
20'b00001101010000000011 : ColourData = 12'hFFF;
20'b00001101100000000011 : ColourData = 12'hFFF;
20'b00001101110000000011 : ColourData = 12'hFFF;
20'b00001110000000000011 : ColourData = 12'hFFF;
20'b00001110010000000011 : ColourData = 12'hFFF;
20'b00001110100000000011 : ColourData = 12'hFFF;
20'b00001110110000000011 : ColourData = 12'hFFF;
20'b00000000000000000100 : ColourData = 12'hFFF;
20'b00000000010000000100 : ColourData = 12'hFFF;
20'b00000000100000000100 : ColourData = 12'hFFF;
20'b00000000110000000100 : ColourData = 12'hFFF;
20'b00000001000000000100 : ColourData = 12'hFFF;
20'b00000001010000000100 : ColourData = 12'hFFF;
20'b00000001100000000100 : ColourData = 12'hFFF;
20'b00000001110000000100 : ColourData = 12'hFFF;
20'b00000010000000000100 : ColourData = 12'hFFF;
20'b00000010010000000100 : ColourData = 12'hFFF;
20'b00000010100000000100 : ColourData = 12'hFFF;
20'b00000010110000000100 : ColourData = 12'hFFF;
20'b00000011000000000100 : ColourData = 12'hFFF;
20'b00000011010000000100 : ColourData = 12'hFFF;
20'b00000011100000000100 : ColourData = 12'hFFF;
20'b00000011110000000100 : ColourData = 12'hFFF;
20'b00000100000000000100 : ColourData = 12'hFFF;
20'b00000100010000000100 : ColourData = 12'hFFF;
20'b00000100100000000100 : ColourData = 12'hFFF;
20'b00000100110000000100 : ColourData = 12'hFFF;
20'b00000101000000000100 : ColourData = 12'hFFF;
20'b00000101010000000100 : ColourData = 12'hFFF;
20'b00000101100000000100 : ColourData = 12'hFFF;
20'b00000101110000000100 : ColourData = 12'hFFF;
20'b00000110000000000100 : ColourData = 12'hFFF;
20'b00000110010000000100 : ColourData = 12'hFFF;
20'b00000110100000000100 : ColourData = 12'hFFF;
20'b00000110110000000100 : ColourData = 12'hAAA;
20'b00000111000000000100 : ColourData = 12'h000;
20'b00000111010000000100 : ColourData = 12'h000;
20'b00000111100000000100 : ColourData = 12'h000;
20'b00000111110000000100 : ColourData = 12'h000;
20'b00001000000000000100 : ColourData = 12'hAAA;
20'b00001000010000000100 : ColourData = 12'hFFF;
20'b00001000100000000100 : ColourData = 12'hFFF;
20'b00001000110000000100 : ColourData = 12'hFFF;
20'b00001001000000000100 : ColourData = 12'hFFF;
20'b00001001010000000100 : ColourData = 12'hFFF;
20'b00001001100000000100 : ColourData = 12'hFFF;
20'b00001001110000000100 : ColourData = 12'hFFF;
20'b00001010000000000100 : ColourData = 12'hFFF;
20'b00001010010000000100 : ColourData = 12'hFFF;
20'b00001010100000000100 : ColourData = 12'hFFF;
20'b00001010110000000100 : ColourData = 12'hFFF;
20'b00001011000000000100 : ColourData = 12'hFFF;
20'b00001011010000000100 : ColourData = 12'hFFF;
20'b00001011100000000100 : ColourData = 12'hFFF;
20'b00001011110000000100 : ColourData = 12'hFFF;
20'b00001100000000000100 : ColourData = 12'hFFF;
20'b00001100010000000100 : ColourData = 12'hFFF;
20'b00001100100000000100 : ColourData = 12'hFFF;
20'b00001100110000000100 : ColourData = 12'hFFF;
20'b00001101000000000100 : ColourData = 12'hFFF;
20'b00001101010000000100 : ColourData = 12'hFFF;
20'b00001101100000000100 : ColourData = 12'hFFF;
20'b00001101110000000100 : ColourData = 12'hFFF;
20'b00001110000000000100 : ColourData = 12'hFFF;
20'b00001110010000000100 : ColourData = 12'hFFF;
20'b00001110100000000100 : ColourData = 12'hFFF;
20'b00001110110000000100 : ColourData = 12'hFFF;
20'b00000000000000000101 : ColourData = 12'hFFF;
20'b00000000010000000101 : ColourData = 12'hFFF;
20'b00000000100000000101 : ColourData = 12'hFFF;
20'b00000000110000000101 : ColourData = 12'hFFF;
20'b00000001000000000101 : ColourData = 12'hFFF;
20'b00000001010000000101 : ColourData = 12'hFFF;
20'b00000001100000000101 : ColourData = 12'hFFF;
20'b00000001110000000101 : ColourData = 12'hFFF;
20'b00000010000000000101 : ColourData = 12'hFFF;
20'b00000010010000000101 : ColourData = 12'hFFF;
20'b00000010100000000101 : ColourData = 12'hFFF;
20'b00000010110000000101 : ColourData = 12'hFFF;
20'b00000011000000000101 : ColourData = 12'hFFF;
20'b00000011010000000101 : ColourData = 12'hFFF;
20'b00000011100000000101 : ColourData = 12'hFFF;
20'b00000011110000000101 : ColourData = 12'hFFF;
20'b00000100000000000101 : ColourData = 12'hFFF;
20'b00000100010000000101 : ColourData = 12'hFFF;
20'b00000100100000000101 : ColourData = 12'hFFF;
20'b00000100110000000101 : ColourData = 12'hFFF;
20'b00000101000000000101 : ColourData = 12'hFFF;
20'b00000101010000000101 : ColourData = 12'hFFF;
20'b00000101100000000101 : ColourData = 12'hFFF;
20'b00000101110000000101 : ColourData = 12'hFFF;
20'b00000110000000000101 : ColourData = 12'hFFF;
20'b00000110010000000101 : ColourData = 12'hFFF;
20'b00000110100000000101 : ColourData = 12'hFFF;
20'b00000110110000000101 : ColourData = 12'hAAA;
20'b00000111000000000101 : ColourData = 12'h000;
20'b00000111010000000101 : ColourData = 12'h000;
20'b00000111100000000101 : ColourData = 12'h000;
20'b00000111110000000101 : ColourData = 12'h000;
20'b00001000000000000101 : ColourData = 12'hAAA;
20'b00001000010000000101 : ColourData = 12'hFFF;
20'b00001000100000000101 : ColourData = 12'hFFF;
20'b00001000110000000101 : ColourData = 12'hFFF;
20'b00001001000000000101 : ColourData = 12'hFFF;
20'b00001001010000000101 : ColourData = 12'hFFF;
20'b00001001100000000101 : ColourData = 12'hFFF;
20'b00001001110000000101 : ColourData = 12'hFFF;
20'b00001010000000000101 : ColourData = 12'hFFF;
20'b00001010010000000101 : ColourData = 12'hFFF;
20'b00001010100000000101 : ColourData = 12'hFFF;
20'b00001010110000000101 : ColourData = 12'hFFF;
20'b00001011000000000101 : ColourData = 12'hFFF;
20'b00001011010000000101 : ColourData = 12'hFFF;
20'b00001011100000000101 : ColourData = 12'hFFF;
20'b00001011110000000101 : ColourData = 12'hFFF;
20'b00001100000000000101 : ColourData = 12'hFFF;
20'b00001100010000000101 : ColourData = 12'hFFF;
20'b00001100100000000101 : ColourData = 12'hFFF;
20'b00001100110000000101 : ColourData = 12'hFFF;
20'b00001101000000000101 : ColourData = 12'hFFF;
20'b00001101010000000101 : ColourData = 12'hFFF;
20'b00001101100000000101 : ColourData = 12'hFFF;
20'b00001101110000000101 : ColourData = 12'hFFF;
20'b00001110000000000101 : ColourData = 12'hFFF;
20'b00001110010000000101 : ColourData = 12'hFFF;
20'b00001110100000000101 : ColourData = 12'hFFF;
20'b00001110110000000101 : ColourData = 12'hFFF;
20'b00000000000000000110 : ColourData = 12'hFFF;
20'b00000000010000000110 : ColourData = 12'hFFF;
20'b00000000100000000110 : ColourData = 12'hFFF;
20'b00000000110000000110 : ColourData = 12'hFFF;
20'b00000001000000000110 : ColourData = 12'hFFF;
20'b00000001010000000110 : ColourData = 12'hFFF;
20'b00000001100000000110 : ColourData = 12'hFFF;
20'b00000001110000000110 : ColourData = 12'hFFF;
20'b00000010000000000110 : ColourData = 12'hFFF;
20'b00000010010000000110 : ColourData = 12'hFFF;
20'b00000010100000000110 : ColourData = 12'hFFF;
20'b00000010110000000110 : ColourData = 12'hFFF;
20'b00000011000000000110 : ColourData = 12'hFFF;
20'b00000011010000000110 : ColourData = 12'hFFF;
20'b00000011100000000110 : ColourData = 12'hFFF;
20'b00000011110000000110 : ColourData = 12'hFFF;
20'b00000100000000000110 : ColourData = 12'hFFF;
20'b00000100010000000110 : ColourData = 12'hFFF;
20'b00000100100000000110 : ColourData = 12'hFFF;
20'b00000100110000000110 : ColourData = 12'hFFF;
20'b00000101000000000110 : ColourData = 12'hFFF;
20'b00000101010000000110 : ColourData = 12'hFFF;
20'b00000101100000000110 : ColourData = 12'hFFF;
20'b00000101110000000110 : ColourData = 12'hFFF;
20'b00000110000000000110 : ColourData = 12'hFFF;
20'b00000110010000000110 : ColourData = 12'hFFF;
20'b00000110100000000110 : ColourData = 12'hFFF;
20'b00000110110000000110 : ColourData = 12'hAAA;
20'b00000111000000000110 : ColourData = 12'h000;
20'b00000111010000000110 : ColourData = 12'h000;
20'b00000111100000000110 : ColourData = 12'h000;
20'b00000111110000000110 : ColourData = 12'h000;
20'b00001000000000000110 : ColourData = 12'hAAA;
20'b00001000010000000110 : ColourData = 12'hFFF;
20'b00001000100000000110 : ColourData = 12'hFFF;
20'b00001000110000000110 : ColourData = 12'hFFF;
20'b00001001000000000110 : ColourData = 12'hFFF;
20'b00001001010000000110 : ColourData = 12'hFFF;
20'b00001001100000000110 : ColourData = 12'hFFF;
20'b00001001110000000110 : ColourData = 12'hFFF;
20'b00001010000000000110 : ColourData = 12'hFFF;
20'b00001010010000000110 : ColourData = 12'hFFF;
20'b00001010100000000110 : ColourData = 12'hFFF;
20'b00001010110000000110 : ColourData = 12'hFFF;
20'b00001011000000000110 : ColourData = 12'hFFF;
20'b00001011010000000110 : ColourData = 12'hFFF;
20'b00001011100000000110 : ColourData = 12'hFFF;
20'b00001011110000000110 : ColourData = 12'hFFF;
20'b00001100000000000110 : ColourData = 12'hFFF;
20'b00001100010000000110 : ColourData = 12'hFFF;
20'b00001100100000000110 : ColourData = 12'hFFF;
20'b00001100110000000110 : ColourData = 12'hFFF;
20'b00001101000000000110 : ColourData = 12'hFFF;
20'b00001101010000000110 : ColourData = 12'hFFF;
20'b00001101100000000110 : ColourData = 12'hFFF;
20'b00001101110000000110 : ColourData = 12'hFFF;
20'b00001110000000000110 : ColourData = 12'hFFF;
20'b00001110010000000110 : ColourData = 12'hFFF;
20'b00001110100000000110 : ColourData = 12'hFFF;
20'b00001110110000000110 : ColourData = 12'hFFF;
20'b00000000000000000111 : ColourData = 12'hFFF;
20'b00000000010000000111 : ColourData = 12'hFFF;
20'b00000000100000000111 : ColourData = 12'hFFF;
20'b00000000110000000111 : ColourData = 12'hFFF;
20'b00000001000000000111 : ColourData = 12'hFFF;
20'b00000001010000000111 : ColourData = 12'hFFF;
20'b00000001100000000111 : ColourData = 12'hFFF;
20'b00000001110000000111 : ColourData = 12'hFFF;
20'b00000010000000000111 : ColourData = 12'hFFF;
20'b00000010010000000111 : ColourData = 12'hFFF;
20'b00000010100000000111 : ColourData = 12'hFFF;
20'b00000010110000000111 : ColourData = 12'hFFF;
20'b00000011000000000111 : ColourData = 12'hFFF;
20'b00000011010000000111 : ColourData = 12'hFFF;
20'b00000011100000000111 : ColourData = 12'hFFF;
20'b00000011110000000111 : ColourData = 12'hFFF;
20'b00000100000000000111 : ColourData = 12'hFFF;
20'b00000100010000000111 : ColourData = 12'hFFF;
20'b00000100100000000111 : ColourData = 12'hFFF;
20'b00000100110000000111 : ColourData = 12'hFFF;
20'b00000101000000000111 : ColourData = 12'hFFF;
20'b00000101010000000111 : ColourData = 12'hFFF;
20'b00000101100000000111 : ColourData = 12'hFFF;
20'b00000101110000000111 : ColourData = 12'hFFF;
20'b00000110000000000111 : ColourData = 12'hFFF;
20'b00000110010000000111 : ColourData = 12'hFFF;
20'b00000110100000000111 : ColourData = 12'hFFF;
20'b00000110110000000111 : ColourData = 12'hAAA;
20'b00000111000000000111 : ColourData = 12'h000;
20'b00000111010000000111 : ColourData = 12'h000;
20'b00000111100000000111 : ColourData = 12'h000;
20'b00000111110000000111 : ColourData = 12'h000;
20'b00001000000000000111 : ColourData = 12'hAAA;
20'b00001000010000000111 : ColourData = 12'hFFF;
20'b00001000100000000111 : ColourData = 12'hFFF;
20'b00001000110000000111 : ColourData = 12'hFFF;
20'b00001001000000000111 : ColourData = 12'hFFF;
20'b00001001010000000111 : ColourData = 12'hFFF;
20'b00001001100000000111 : ColourData = 12'hFFF;
20'b00001001110000000111 : ColourData = 12'hFFF;
20'b00001010000000000111 : ColourData = 12'hFFF;
20'b00001010010000000111 : ColourData = 12'hFFF;
20'b00001010100000000111 : ColourData = 12'hFFF;
20'b00001010110000000111 : ColourData = 12'hFFF;
20'b00001011000000000111 : ColourData = 12'hFFF;
20'b00001011010000000111 : ColourData = 12'hFFF;
20'b00001011100000000111 : ColourData = 12'hFFF;
20'b00001011110000000111 : ColourData = 12'hFFF;
20'b00001100000000000111 : ColourData = 12'hFFF;
20'b00001100010000000111 : ColourData = 12'hFFF;
20'b00001100100000000111 : ColourData = 12'hFFF;
20'b00001100110000000111 : ColourData = 12'hFFF;
20'b00001101000000000111 : ColourData = 12'hFFF;
20'b00001101010000000111 : ColourData = 12'hFFF;
20'b00001101100000000111 : ColourData = 12'hFFF;
20'b00001101110000000111 : ColourData = 12'hFFF;
20'b00001110000000000111 : ColourData = 12'hFFF;
20'b00001110010000000111 : ColourData = 12'hFFF;
20'b00001110100000000111 : ColourData = 12'hFFF;
20'b00001110110000000111 : ColourData = 12'hFFF;
20'b00000000000000001000 : ColourData = 12'hFFF;
20'b00000000010000001000 : ColourData = 12'hFFF;
20'b00000000100000001000 : ColourData = 12'hFFF;
20'b00000000110000001000 : ColourData = 12'hFFF;
20'b00000001000000001000 : ColourData = 12'hFFF;
20'b00000001010000001000 : ColourData = 12'hFFF;
20'b00000001100000001000 : ColourData = 12'hFFF;
20'b00000001110000001000 : ColourData = 12'hFFF;
20'b00000010000000001000 : ColourData = 12'hFFF;
20'b00000010010000001000 : ColourData = 12'hFFF;
20'b00000010100000001000 : ColourData = 12'hFFF;
20'b00000010110000001000 : ColourData = 12'hFFF;
20'b00000011000000001000 : ColourData = 12'hFFF;
20'b00000011010000001000 : ColourData = 12'hFFF;
20'b00000011100000001000 : ColourData = 12'hFFF;
20'b00000011110000001000 : ColourData = 12'hFFF;
20'b00000100000000001000 : ColourData = 12'hFFF;
20'b00000100010000001000 : ColourData = 12'hFFF;
20'b00000100100000001000 : ColourData = 12'hFFF;
20'b00000100110000001000 : ColourData = 12'hFFF;
20'b00000101000000001000 : ColourData = 12'hFFF;
20'b00000101010000001000 : ColourData = 12'hFFF;
20'b00000101100000001000 : ColourData = 12'hFFF;
20'b00000101110000001000 : ColourData = 12'hFFF;
20'b00000110000000001000 : ColourData = 12'hFFF;
20'b00000110010000001000 : ColourData = 12'hFFF;
20'b00000110100000001000 : ColourData = 12'hFFF;
20'b00000110110000001000 : ColourData = 12'hAAA;
20'b00000111000000001000 : ColourData = 12'h000;
20'b00000111010000001000 : ColourData = 12'h000;
20'b00000111100000001000 : ColourData = 12'h000;
20'b00000111110000001000 : ColourData = 12'h000;
20'b00001000000000001000 : ColourData = 12'hAAA;
20'b00001000010000001000 : ColourData = 12'hFFF;
20'b00001000100000001000 : ColourData = 12'hFFF;
20'b00001000110000001000 : ColourData = 12'hFFF;
20'b00001001000000001000 : ColourData = 12'hFFF;
20'b00001001010000001000 : ColourData = 12'hFFF;
20'b00001001100000001000 : ColourData = 12'hFFF;
20'b00001001110000001000 : ColourData = 12'hFFF;
20'b00001010000000001000 : ColourData = 12'hFFF;
20'b00001010010000001000 : ColourData = 12'hFFF;
20'b00001010100000001000 : ColourData = 12'hFFF;
20'b00001010110000001000 : ColourData = 12'hFFF;
20'b00001011000000001000 : ColourData = 12'hFFF;
20'b00001011010000001000 : ColourData = 12'hFFF;
20'b00001011100000001000 : ColourData = 12'hFFF;
20'b00001011110000001000 : ColourData = 12'hFFF;
20'b00001100000000001000 : ColourData = 12'hFFF;
20'b00001100010000001000 : ColourData = 12'hFFF;
20'b00001100100000001000 : ColourData = 12'hFFF;
20'b00001100110000001000 : ColourData = 12'hFFF;
20'b00001101000000001000 : ColourData = 12'hFFF;
20'b00001101010000001000 : ColourData = 12'hFFF;
20'b00001101100000001000 : ColourData = 12'hFFF;
20'b00001101110000001000 : ColourData = 12'hFFF;
20'b00001110000000001000 : ColourData = 12'hFFF;
20'b00001110010000001000 : ColourData = 12'hFFF;
20'b00001110100000001000 : ColourData = 12'hFFF;
20'b00001110110000001000 : ColourData = 12'hFFF;
20'b00000000000000001001 : ColourData = 12'hFFF;
20'b00000000010000001001 : ColourData = 12'hFFF;
20'b00000000100000001001 : ColourData = 12'hFFF;
20'b00000000110000001001 : ColourData = 12'hFFF;
20'b00000001000000001001 : ColourData = 12'hFFF;
20'b00000001010000001001 : ColourData = 12'hFFF;
20'b00000001100000001001 : ColourData = 12'hFFF;
20'b00000001110000001001 : ColourData = 12'hFFF;
20'b00000010000000001001 : ColourData = 12'hFFF;
20'b00000010010000001001 : ColourData = 12'hFFF;
20'b00000010100000001001 : ColourData = 12'hFFF;
20'b00000010110000001001 : ColourData = 12'hFFF;
20'b00000011000000001001 : ColourData = 12'hFFF;
20'b00000011010000001001 : ColourData = 12'hFFF;
20'b00000011100000001001 : ColourData = 12'hFFF;
20'b00000011110000001001 : ColourData = 12'hFFF;
20'b00000100000000001001 : ColourData = 12'hFFF;
20'b00000100010000001001 : ColourData = 12'hFFF;
20'b00000100100000001001 : ColourData = 12'hFFF;
20'b00000100110000001001 : ColourData = 12'hFFF;
20'b00000101000000001001 : ColourData = 12'hFFF;
20'b00000101010000001001 : ColourData = 12'hFFF;
20'b00000101100000001001 : ColourData = 12'hFFF;
20'b00000101110000001001 : ColourData = 12'hFFF;
20'b00000110000000001001 : ColourData = 12'hFFF;
20'b00000110010000001001 : ColourData = 12'hFFF;
20'b00000110100000001001 : ColourData = 12'hFFF;
20'b00000110110000001001 : ColourData = 12'hAAA;
20'b00000111000000001001 : ColourData = 12'h000;
20'b00000111010000001001 : ColourData = 12'h000;
20'b00000111100000001001 : ColourData = 12'h000;
20'b00000111110000001001 : ColourData = 12'h000;
20'b00001000000000001001 : ColourData = 12'hAAA;
20'b00001000010000001001 : ColourData = 12'hFFF;
20'b00001000100000001001 : ColourData = 12'hFFF;
20'b00001000110000001001 : ColourData = 12'hFFF;
20'b00001001000000001001 : ColourData = 12'hFFF;
20'b00001001010000001001 : ColourData = 12'hFFF;
20'b00001001100000001001 : ColourData = 12'hFFF;
20'b00001001110000001001 : ColourData = 12'hFFF;
20'b00001010000000001001 : ColourData = 12'hFFF;
20'b00001010010000001001 : ColourData = 12'hFFF;
20'b00001010100000001001 : ColourData = 12'hFFF;
20'b00001010110000001001 : ColourData = 12'hFFF;
20'b00001011000000001001 : ColourData = 12'hFFF;
20'b00001011010000001001 : ColourData = 12'hFFF;
20'b00001011100000001001 : ColourData = 12'hFFF;
20'b00001011110000001001 : ColourData = 12'hFFF;
20'b00001100000000001001 : ColourData = 12'hFFF;
20'b00001100010000001001 : ColourData = 12'hFFF;
20'b00001100100000001001 : ColourData = 12'hFFF;
20'b00001100110000001001 : ColourData = 12'hFFF;
20'b00001101000000001001 : ColourData = 12'hFFF;
20'b00001101010000001001 : ColourData = 12'hFFF;
20'b00001101100000001001 : ColourData = 12'hFFF;
20'b00001101110000001001 : ColourData = 12'hFFF;
20'b00001110000000001001 : ColourData = 12'hFFF;
20'b00001110010000001001 : ColourData = 12'hFFF;
20'b00001110100000001001 : ColourData = 12'hFFF;
20'b00001110110000001001 : ColourData = 12'hFFF;
20'b00000000000000001010 : ColourData = 12'hFFF;
20'b00000000010000001010 : ColourData = 12'hFFF;
20'b00000000100000001010 : ColourData = 12'hFFF;
20'b00000000110000001010 : ColourData = 12'hFFF;
20'b00000001000000001010 : ColourData = 12'hFFF;
20'b00000001010000001010 : ColourData = 12'hFFF;
20'b00000001100000001010 : ColourData = 12'hFFF;
20'b00000001110000001010 : ColourData = 12'hFFF;
20'b00000010000000001010 : ColourData = 12'hFFF;
20'b00000010010000001010 : ColourData = 12'hFFF;
20'b00000010100000001010 : ColourData = 12'hFFF;
20'b00000010110000001010 : ColourData = 12'hFFF;
20'b00000011000000001010 : ColourData = 12'hFFF;
20'b00000011010000001010 : ColourData = 12'hFFF;
20'b00000011100000001010 : ColourData = 12'hFFF;
20'b00000011110000001010 : ColourData = 12'hFFF;
20'b00000100000000001010 : ColourData = 12'hFFF;
20'b00000100010000001010 : ColourData = 12'hFFF;
20'b00000100100000001010 : ColourData = 12'hDEC;
20'b00000100110000001010 : ColourData = 12'hBD9;
20'b00000101000000001010 : ColourData = 12'hBD9;
20'b00000101010000001010 : ColourData = 12'hBD9;
20'b00000101100000001010 : ColourData = 12'hBD9;
20'b00000101110000001010 : ColourData = 12'hBD9;
20'b00000110000000001010 : ColourData = 12'hBD9;
20'b00000110010000001010 : ColourData = 12'hBD9;
20'b00000110100000001010 : ColourData = 12'hCEA;
20'b00000110110000001010 : ColourData = 12'h896;
20'b00000111000000001010 : ColourData = 12'h000;
20'b00000111010000001010 : ColourData = 12'h000;
20'b00000111100000001010 : ColourData = 12'h000;
20'b00000111110000001010 : ColourData = 12'h000;
20'b00001000000000001010 : ColourData = 12'h896;
20'b00001000010000001010 : ColourData = 12'hCEA;
20'b00001000100000001010 : ColourData = 12'hBD9;
20'b00001000110000001010 : ColourData = 12'hBD9;
20'b00001001000000001010 : ColourData = 12'hBD9;
20'b00001001010000001010 : ColourData = 12'hBD9;
20'b00001001100000001010 : ColourData = 12'hBD9;
20'b00001001110000001010 : ColourData = 12'hBD9;
20'b00001010000000001010 : ColourData = 12'hBD9;
20'b00001010010000001010 : ColourData = 12'hDEC;
20'b00001010100000001010 : ColourData = 12'hFFF;
20'b00001010110000001010 : ColourData = 12'hFFF;
20'b00001011000000001010 : ColourData = 12'hFFF;
20'b00001011010000001010 : ColourData = 12'hFFF;
20'b00001011100000001010 : ColourData = 12'hFFF;
20'b00001011110000001010 : ColourData = 12'hFFF;
20'b00001100000000001010 : ColourData = 12'hFFF;
20'b00001100010000001010 : ColourData = 12'hFFF;
20'b00001100100000001010 : ColourData = 12'hFFF;
20'b00001100110000001010 : ColourData = 12'hFFF;
20'b00001101000000001010 : ColourData = 12'hFFF;
20'b00001101010000001010 : ColourData = 12'hFFF;
20'b00001101100000001010 : ColourData = 12'hFFF;
20'b00001101110000001010 : ColourData = 12'hFFF;
20'b00001110000000001010 : ColourData = 12'hFFF;
20'b00001110010000001010 : ColourData = 12'hFFF;
20'b00001110100000001010 : ColourData = 12'hFFF;
20'b00001110110000001010 : ColourData = 12'hFFF;
20'b00000000000000001011 : ColourData = 12'hFFF;
20'b00000000010000001011 : ColourData = 12'hFFF;
20'b00000000100000001011 : ColourData = 12'hFFF;
20'b00000000110000001011 : ColourData = 12'hFFF;
20'b00000001000000001011 : ColourData = 12'hFFF;
20'b00000001010000001011 : ColourData = 12'hFFF;
20'b00000001100000001011 : ColourData = 12'hFFF;
20'b00000001110000001011 : ColourData = 12'hFFF;
20'b00000010000000001011 : ColourData = 12'hFFF;
20'b00000010010000001011 : ColourData = 12'hFFF;
20'b00000010100000001011 : ColourData = 12'hFFF;
20'b00000010110000001011 : ColourData = 12'hFFF;
20'b00000011000000001011 : ColourData = 12'hFFF;
20'b00000011010000001011 : ColourData = 12'hFFF;
20'b00000011100000001011 : ColourData = 12'hFFF;
20'b00000011110000001011 : ColourData = 12'hFFF;
20'b00000100000000001011 : ColourData = 12'hFFF;
20'b00000100010000001011 : ColourData = 12'hFFF;
20'b00000100100000001011 : ColourData = 12'h9C7;
20'b00000100110000001011 : ColourData = 12'h490;
20'b00000101000000001011 : ColourData = 12'h590;
20'b00000101010000001011 : ColourData = 12'h590;
20'b00000101100000001011 : ColourData = 12'h590;
20'b00000101110000001011 : ColourData = 12'h590;
20'b00000110000000001011 : ColourData = 12'h590;
20'b00000110010000001011 : ColourData = 12'h590;
20'b00000110100000001011 : ColourData = 12'h5A0;
20'b00000110110000001011 : ColourData = 12'h360;
20'b00000111000000001011 : ColourData = 12'h000;
20'b00000111010000001011 : ColourData = 12'h000;
20'b00000111100000001011 : ColourData = 12'h000;
20'b00000111110000001011 : ColourData = 12'h000;
20'b00001000000000001011 : ColourData = 12'h360;
20'b00001000010000001011 : ColourData = 12'h5A0;
20'b00001000100000001011 : ColourData = 12'h590;
20'b00001000110000001011 : ColourData = 12'h590;
20'b00001001000000001011 : ColourData = 12'h590;
20'b00001001010000001011 : ColourData = 12'h590;
20'b00001001100000001011 : ColourData = 12'h590;
20'b00001001110000001011 : ColourData = 12'h590;
20'b00001010000000001011 : ColourData = 12'h490;
20'b00001010010000001011 : ColourData = 12'h9C7;
20'b00001010100000001011 : ColourData = 12'hFFF;
20'b00001010110000001011 : ColourData = 12'hFFF;
20'b00001011000000001011 : ColourData = 12'hFFF;
20'b00001011010000001011 : ColourData = 12'hFFF;
20'b00001011100000001011 : ColourData = 12'hFFF;
20'b00001011110000001011 : ColourData = 12'hFFF;
20'b00001100000000001011 : ColourData = 12'hFFF;
20'b00001100010000001011 : ColourData = 12'hFFF;
20'b00001100100000001011 : ColourData = 12'hFFF;
20'b00001100110000001011 : ColourData = 12'hFFF;
20'b00001101000000001011 : ColourData = 12'hFFF;
20'b00001101010000001011 : ColourData = 12'hFFF;
20'b00001101100000001011 : ColourData = 12'hFFF;
20'b00001101110000001011 : ColourData = 12'hFFF;
20'b00001110000000001011 : ColourData = 12'hFFF;
20'b00001110010000001011 : ColourData = 12'hFFF;
20'b00001110100000001011 : ColourData = 12'hFFF;
20'b00001110110000001011 : ColourData = 12'hFFF;
20'b00000000000000001100 : ColourData = 12'hFFF;
20'b00000000010000001100 : ColourData = 12'hFFF;
20'b00000000100000001100 : ColourData = 12'hFFF;
20'b00000000110000001100 : ColourData = 12'hFFF;
20'b00000001000000001100 : ColourData = 12'hFFF;
20'b00000001010000001100 : ColourData = 12'hFFF;
20'b00000001100000001100 : ColourData = 12'hFFF;
20'b00000001110000001100 : ColourData = 12'hFFF;
20'b00000010000000001100 : ColourData = 12'hFFF;
20'b00000010010000001100 : ColourData = 12'hFFF;
20'b00000010100000001100 : ColourData = 12'hFFF;
20'b00000010110000001100 : ColourData = 12'hFFF;
20'b00000011000000001100 : ColourData = 12'hFFF;
20'b00000011010000001100 : ColourData = 12'hEEE;
20'b00000011100000001100 : ColourData = 12'h8B5;
20'b00000011110000001100 : ColourData = 12'h8B6;
20'b00000100000000001100 : ColourData = 12'h8B6;
20'b00000100010000001100 : ColourData = 12'h9B6;
20'b00000100100000001100 : ColourData = 12'h7A3;
20'b00000100110000001100 : ColourData = 12'h591;
20'b00000101000000001100 : ColourData = 12'h5A1;
20'b00000101010000001100 : ColourData = 12'h5A1;
20'b00000101100000001100 : ColourData = 12'h5A1;
20'b00000101110000001100 : ColourData = 12'h5A1;
20'b00000110000000001100 : ColourData = 12'h5A1;
20'b00000110010000001100 : ColourData = 12'h5A1;
20'b00000110100000001100 : ColourData = 12'h6A1;
20'b00000110110000001100 : ColourData = 12'h360;
20'b00000111000000001100 : ColourData = 12'h000;
20'b00000111010000001100 : ColourData = 12'h000;
20'b00000111100000001100 : ColourData = 12'h000;
20'b00000111110000001100 : ColourData = 12'h000;
20'b00001000000000001100 : ColourData = 12'h360;
20'b00001000010000001100 : ColourData = 12'h6A1;
20'b00001000100000001100 : ColourData = 12'h5A1;
20'b00001000110000001100 : ColourData = 12'h5A1;
20'b00001001000000001100 : ColourData = 12'h5A1;
20'b00001001010000001100 : ColourData = 12'h5A1;
20'b00001001100000001100 : ColourData = 12'h5A1;
20'b00001001110000001100 : ColourData = 12'h5A1;
20'b00001010000000001100 : ColourData = 12'h591;
20'b00001010010000001100 : ColourData = 12'h7A3;
20'b00001010100000001100 : ColourData = 12'h9B6;
20'b00001010110000001100 : ColourData = 12'h8B6;
20'b00001011000000001100 : ColourData = 12'h8B6;
20'b00001011010000001100 : ColourData = 12'h8B5;
20'b00001011100000001100 : ColourData = 12'hEEE;
20'b00001011110000001100 : ColourData = 12'hFFF;
20'b00001100000000001100 : ColourData = 12'hFFF;
20'b00001100010000001100 : ColourData = 12'hFFF;
20'b00001100100000001100 : ColourData = 12'hFFF;
20'b00001100110000001100 : ColourData = 12'hFFF;
20'b00001101000000001100 : ColourData = 12'hFFF;
20'b00001101010000001100 : ColourData = 12'hFFF;
20'b00001101100000001100 : ColourData = 12'hFFF;
20'b00001101110000001100 : ColourData = 12'hFFF;
20'b00001110000000001100 : ColourData = 12'hFFF;
20'b00001110010000001100 : ColourData = 12'hFFF;
20'b00001110100000001100 : ColourData = 12'hFFF;
20'b00001110110000001100 : ColourData = 12'hFFF;
20'b00000000000000001101 : ColourData = 12'hFFF;
20'b00000000010000001101 : ColourData = 12'hFFF;
20'b00000000100000001101 : ColourData = 12'hFFF;
20'b00000000110000001101 : ColourData = 12'hFFF;
20'b00000001000000001101 : ColourData = 12'hFFF;
20'b00000001010000001101 : ColourData = 12'hFFF;
20'b00000001100000001101 : ColourData = 12'hFFF;
20'b00000001110000001101 : ColourData = 12'hFFF;
20'b00000010000000001101 : ColourData = 12'hFFF;
20'b00000010010000001101 : ColourData = 12'hFFF;
20'b00000010100000001101 : ColourData = 12'hFFF;
20'b00000010110000001101 : ColourData = 12'hFFF;
20'b00000011000000001101 : ColourData = 12'hFFF;
20'b00000011010000001101 : ColourData = 12'hDED;
20'b00000011100000001101 : ColourData = 12'h590;
20'b00000011110000001101 : ColourData = 12'h590;
20'b00000100000000001101 : ColourData = 12'h590;
20'b00000100010000001101 : ColourData = 12'h590;
20'b00000100100000001101 : ColourData = 12'h5A1;
20'b00000100110000001101 : ColourData = 12'h5A1;
20'b00000101000000001101 : ColourData = 12'h5A1;
20'b00000101010000001101 : ColourData = 12'h5A1;
20'b00000101100000001101 : ColourData = 12'h5A1;
20'b00000101110000001101 : ColourData = 12'h5A1;
20'b00000110000000001101 : ColourData = 12'h5A1;
20'b00000110010000001101 : ColourData = 12'h5A1;
20'b00000110100000001101 : ColourData = 12'h6A1;
20'b00000110110000001101 : ColourData = 12'h360;
20'b00000111000000001101 : ColourData = 12'h000;
20'b00000111010000001101 : ColourData = 12'h000;
20'b00000111100000001101 : ColourData = 12'h000;
20'b00000111110000001101 : ColourData = 12'h000;
20'b00001000000000001101 : ColourData = 12'h360;
20'b00001000010000001101 : ColourData = 12'h6A1;
20'b00001000100000001101 : ColourData = 12'h5A1;
20'b00001000110000001101 : ColourData = 12'h5A1;
20'b00001001000000001101 : ColourData = 12'h5A1;
20'b00001001010000001101 : ColourData = 12'h5A1;
20'b00001001100000001101 : ColourData = 12'h5A1;
20'b00001001110000001101 : ColourData = 12'h5A1;
20'b00001010000000001101 : ColourData = 12'h5A1;
20'b00001010010000001101 : ColourData = 12'h5A1;
20'b00001010100000001101 : ColourData = 12'h590;
20'b00001010110000001101 : ColourData = 12'h590;
20'b00001011000000001101 : ColourData = 12'h590;
20'b00001011010000001101 : ColourData = 12'h590;
20'b00001011100000001101 : ColourData = 12'hDED;
20'b00001011110000001101 : ColourData = 12'hFFF;
20'b00001100000000001101 : ColourData = 12'hFFF;
20'b00001100010000001101 : ColourData = 12'hFFF;
20'b00001100100000001101 : ColourData = 12'hFFF;
20'b00001100110000001101 : ColourData = 12'hFFF;
20'b00001101000000001101 : ColourData = 12'hFFF;
20'b00001101010000001101 : ColourData = 12'hFFF;
20'b00001101100000001101 : ColourData = 12'hFFF;
20'b00001101110000001101 : ColourData = 12'hFFF;
20'b00001110000000001101 : ColourData = 12'hFFF;
20'b00001110010000001101 : ColourData = 12'hFFF;
20'b00001110100000001101 : ColourData = 12'hFFF;
20'b00001110110000001101 : ColourData = 12'hFFF;
20'b00000000000000001110 : ColourData = 12'hFFF;
20'b00000000010000001110 : ColourData = 12'hFFF;
20'b00000000100000001110 : ColourData = 12'hFFF;
20'b00000000110000001110 : ColourData = 12'hFFF;
20'b00000001000000001110 : ColourData = 12'hBBB;
20'b00000001010000001110 : ColourData = 12'h444;
20'b00000001100000001110 : ColourData = 12'h555;
20'b00000001110000001110 : ColourData = 12'h555;
20'b00000010000000001110 : ColourData = 12'h555;
20'b00000010010000001110 : ColourData = 12'h555;
20'b00000010100000001110 : ColourData = 12'h555;
20'b00000010110000001110 : ColourData = 12'h555;
20'b00000011000000001110 : ColourData = 12'h555;
20'b00000011010000001110 : ColourData = 12'h454;
20'b00000011100000001110 : ColourData = 12'h360;
20'b00000011110000001110 : ColourData = 12'h360;
20'b00000100000000001110 : ColourData = 12'h360;
20'b00000100010000001110 : ColourData = 12'h360;
20'b00000100100000001110 : ColourData = 12'h360;
20'b00000100110000001110 : ColourData = 12'h360;
20'b00000101000000001110 : ColourData = 12'h360;
20'b00000101010000001110 : ColourData = 12'h360;
20'b00000101100000001110 : ColourData = 12'h360;
20'b00000101110000001110 : ColourData = 12'h360;
20'b00000110000000001110 : ColourData = 12'h360;
20'b00000110010000001110 : ColourData = 12'h360;
20'b00000110100000001110 : ColourData = 12'h470;
20'b00000110110000001110 : ColourData = 12'h240;
20'b00000111000000001110 : ColourData = 12'h000;
20'b00000111010000001110 : ColourData = 12'h000;
20'b00000111100000001110 : ColourData = 12'h000;
20'b00000111110000001110 : ColourData = 12'h000;
20'b00001000000000001110 : ColourData = 12'h240;
20'b00001000010000001110 : ColourData = 12'h470;
20'b00001000100000001110 : ColourData = 12'h360;
20'b00001000110000001110 : ColourData = 12'h360;
20'b00001001000000001110 : ColourData = 12'h360;
20'b00001001010000001110 : ColourData = 12'h360;
20'b00001001100000001110 : ColourData = 12'h360;
20'b00001001110000001110 : ColourData = 12'h360;
20'b00001010000000001110 : ColourData = 12'h360;
20'b00001010010000001110 : ColourData = 12'h360;
20'b00001010100000001110 : ColourData = 12'h360;
20'b00001010110000001110 : ColourData = 12'h360;
20'b00001011000000001110 : ColourData = 12'h360;
20'b00001011010000001110 : ColourData = 12'h360;
20'b00001011100000001110 : ColourData = 12'h454;
20'b00001011110000001110 : ColourData = 12'h555;
20'b00001100000000001110 : ColourData = 12'h555;
20'b00001100010000001110 : ColourData = 12'h555;
20'b00001100100000001110 : ColourData = 12'h555;
20'b00001100110000001110 : ColourData = 12'h555;
20'b00001101000000001110 : ColourData = 12'h555;
20'b00001101010000001110 : ColourData = 12'h555;
20'b00001101100000001110 : ColourData = 12'h444;
20'b00001101110000001110 : ColourData = 12'hBBB;
20'b00001110000000001110 : ColourData = 12'hFFF;
20'b00001110010000001110 : ColourData = 12'hFFF;
20'b00001110100000001110 : ColourData = 12'hFFF;
20'b00001110110000001110 : ColourData = 12'hFFF;
20'b00000000000000001111 : ColourData = 12'hFFF;
20'b00000000010000001111 : ColourData = 12'hFFF;
20'b00000000100000001111 : ColourData = 12'hFFF;
20'b00000000110000001111 : ColourData = 12'hFFF;
20'b00000001000000001111 : ColourData = 12'hAAA;
20'b00000001010000001111 : ColourData = 12'h222;
20'b00000001100000001111 : ColourData = 12'h333;
20'b00000001110000001111 : ColourData = 12'h333;
20'b00000010000000001111 : ColourData = 12'h333;
20'b00000010010000001111 : ColourData = 12'h333;
20'b00000010100000001111 : ColourData = 12'h333;
20'b00000010110000001111 : ColourData = 12'h333;
20'b00000011000000001111 : ColourData = 12'h333;
20'b00000011010000001111 : ColourData = 12'h333;
20'b00000011100000001111 : ColourData = 12'h360;
20'b00000011110000001111 : ColourData = 12'h360;
20'b00000100000000001111 : ColourData = 12'h360;
20'b00000100010000001111 : ColourData = 12'h360;
20'b00000100100000001111 : ColourData = 12'h360;
20'b00000100110000001111 : ColourData = 12'h360;
20'b00000101000000001111 : ColourData = 12'h360;
20'b00000101010000001111 : ColourData = 12'h360;
20'b00000101100000001111 : ColourData = 12'h360;
20'b00000101110000001111 : ColourData = 12'h360;
20'b00000110000000001111 : ColourData = 12'h360;
20'b00000110010000001111 : ColourData = 12'h360;
20'b00000110100000001111 : ColourData = 12'h360;
20'b00000110110000001111 : ColourData = 12'h240;
20'b00000111000000001111 : ColourData = 12'h000;
20'b00000111010000001111 : ColourData = 12'h000;
20'b00000111100000001111 : ColourData = 12'h000;
20'b00000111110000001111 : ColourData = 12'h000;
20'b00001000000000001111 : ColourData = 12'h240;
20'b00001000010000001111 : ColourData = 12'h360;
20'b00001000100000001111 : ColourData = 12'h360;
20'b00001000110000001111 : ColourData = 12'h360;
20'b00001001000000001111 : ColourData = 12'h360;
20'b00001001010000001111 : ColourData = 12'h360;
20'b00001001100000001111 : ColourData = 12'h360;
20'b00001001110000001111 : ColourData = 12'h360;
20'b00001010000000001111 : ColourData = 12'h360;
20'b00001010010000001111 : ColourData = 12'h360;
20'b00001010100000001111 : ColourData = 12'h360;
20'b00001010110000001111 : ColourData = 12'h360;
20'b00001011000000001111 : ColourData = 12'h360;
20'b00001011010000001111 : ColourData = 12'h360;
20'b00001011100000001111 : ColourData = 12'h333;
20'b00001011110000001111 : ColourData = 12'h333;
20'b00001100000000001111 : ColourData = 12'h333;
20'b00001100010000001111 : ColourData = 12'h333;
20'b00001100100000001111 : ColourData = 12'h333;
20'b00001100110000001111 : ColourData = 12'h333;
20'b00001101000000001111 : ColourData = 12'h333;
20'b00001101010000001111 : ColourData = 12'h333;
20'b00001101100000001111 : ColourData = 12'h222;
20'b00001101110000001111 : ColourData = 12'hAAA;
20'b00001110000000001111 : ColourData = 12'hFFF;
20'b00001110010000001111 : ColourData = 12'hFFF;
20'b00001110100000001111 : ColourData = 12'hFFF;
20'b00001110110000001111 : ColourData = 12'hFFF;
20'b00000000000000010000 : ColourData = 12'hFFF;
20'b00000000010000010000 : ColourData = 12'hFFF;
20'b00000000100000010000 : ColourData = 12'hFFF;
20'b00000000110000010000 : ColourData = 12'hFFF;
20'b00000001000000010000 : ColourData = 12'h999;
20'b00000001010000010000 : ColourData = 12'h000;
20'b00000001100000010000 : ColourData = 12'h000;
20'b00000001110000010000 : ColourData = 12'h000;
20'b00000010000000010000 : ColourData = 12'h000;
20'b00000010010000010000 : ColourData = 12'h000;
20'b00000010100000010000 : ColourData = 12'h000;
20'b00000010110000010000 : ColourData = 12'h000;
20'b00000011000000010000 : ColourData = 12'h000;
20'b00000011010000010000 : ColourData = 12'h000;
20'b00000011100000010000 : ColourData = 12'h360;
20'b00000011110000010000 : ColourData = 12'h360;
20'b00000100000000010000 : ColourData = 12'h360;
20'b00000100010000010000 : ColourData = 12'h360;
20'b00000100100000010000 : ColourData = 12'h360;
20'b00000100110000010000 : ColourData = 12'h360;
20'b00000101000000010000 : ColourData = 12'h360;
20'b00000101010000010000 : ColourData = 12'h360;
20'b00000101100000010000 : ColourData = 12'h360;
20'b00000101110000010000 : ColourData = 12'h360;
20'b00000110000000010000 : ColourData = 12'h360;
20'b00000110010000010000 : ColourData = 12'h360;
20'b00000110100000010000 : ColourData = 12'h360;
20'b00000110110000010000 : ColourData = 12'h240;
20'b00000111000000010000 : ColourData = 12'h000;
20'b00000111010000010000 : ColourData = 12'h000;
20'b00000111100000010000 : ColourData = 12'h000;
20'b00000111110000010000 : ColourData = 12'h000;
20'b00001000000000010000 : ColourData = 12'h240;
20'b00001000010000010000 : ColourData = 12'h360;
20'b00001000100000010000 : ColourData = 12'h360;
20'b00001000110000010000 : ColourData = 12'h360;
20'b00001001000000010000 : ColourData = 12'h360;
20'b00001001010000010000 : ColourData = 12'h360;
20'b00001001100000010000 : ColourData = 12'h360;
20'b00001001110000010000 : ColourData = 12'h360;
20'b00001010000000010000 : ColourData = 12'h360;
20'b00001010010000010000 : ColourData = 12'h360;
20'b00001010100000010000 : ColourData = 12'h360;
20'b00001010110000010000 : ColourData = 12'h360;
20'b00001011000000010000 : ColourData = 12'h360;
20'b00001011010000010000 : ColourData = 12'h360;
20'b00001011100000010000 : ColourData = 12'h000;
20'b00001011110000010000 : ColourData = 12'h000;
20'b00001100000000010000 : ColourData = 12'h000;
20'b00001100010000010000 : ColourData = 12'h000;
20'b00001100100000010000 : ColourData = 12'h000;
20'b00001100110000010000 : ColourData = 12'h000;
20'b00001101000000010000 : ColourData = 12'h000;
20'b00001101010000010000 : ColourData = 12'h000;
20'b00001101100000010000 : ColourData = 12'h000;
20'b00001101110000010000 : ColourData = 12'h999;
20'b00001110000000010000 : ColourData = 12'hFFF;
20'b00001110010000010000 : ColourData = 12'hFFF;
20'b00001110100000010000 : ColourData = 12'hFFF;
20'b00001110110000010000 : ColourData = 12'hFFF;
20'b00000000000000010001 : ColourData = 12'hBBB;
20'b00000000010000010001 : ColourData = 12'hBBB;
20'b00000000100000010001 : ColourData = 12'hBBB;
20'b00000000110000010001 : ColourData = 12'hCCC;
20'b00000001000000010001 : ColourData = 12'h777;
20'b00000001010000010001 : ColourData = 12'h000;
20'b00000001100000010001 : ColourData = 12'h000;
20'b00000001110000010001 : ColourData = 12'h000;
20'b00000010000000010001 : ColourData = 12'h000;
20'b00000010010000010001 : ColourData = 12'h000;
20'b00000010100000010001 : ColourData = 12'h000;
20'b00000010110000010001 : ColourData = 12'h000;
20'b00000011000000010001 : ColourData = 12'h000;
20'b00000011010000010001 : ColourData = 12'h110;
20'b00000011100000010001 : ColourData = 12'h360;
20'b00000011110000010001 : ColourData = 12'h360;
20'b00000100000000010001 : ColourData = 12'h360;
20'b00000100010000010001 : ColourData = 12'h360;
20'b00000100100000010001 : ColourData = 12'h360;
20'b00000100110000010001 : ColourData = 12'h360;
20'b00000101000000010001 : ColourData = 12'h360;
20'b00000101010000010001 : ColourData = 12'h360;
20'b00000101100000010001 : ColourData = 12'h360;
20'b00000101110000010001 : ColourData = 12'h360;
20'b00000110000000010001 : ColourData = 12'h360;
20'b00000110010000010001 : ColourData = 12'h360;
20'b00000110100000010001 : ColourData = 12'h360;
20'b00000110110000010001 : ColourData = 12'h240;
20'b00000111000000010001 : ColourData = 12'h000;
20'b00000111010000010001 : ColourData = 12'h000;
20'b00000111100000010001 : ColourData = 12'h000;
20'b00000111110000010001 : ColourData = 12'h000;
20'b00001000000000010001 : ColourData = 12'h240;
20'b00001000010000010001 : ColourData = 12'h360;
20'b00001000100000010001 : ColourData = 12'h360;
20'b00001000110000010001 : ColourData = 12'h360;
20'b00001001000000010001 : ColourData = 12'h360;
20'b00001001010000010001 : ColourData = 12'h360;
20'b00001001100000010001 : ColourData = 12'h360;
20'b00001001110000010001 : ColourData = 12'h360;
20'b00001010000000010001 : ColourData = 12'h360;
20'b00001010010000010001 : ColourData = 12'h360;
20'b00001010100000010001 : ColourData = 12'h360;
20'b00001010110000010001 : ColourData = 12'h360;
20'b00001011000000010001 : ColourData = 12'h360;
20'b00001011010000010001 : ColourData = 12'h360;
20'b00001011100000010001 : ColourData = 12'h110;
20'b00001011110000010001 : ColourData = 12'h000;
20'b00001100000000010001 : ColourData = 12'h000;
20'b00001100010000010001 : ColourData = 12'h000;
20'b00001100100000010001 : ColourData = 12'h000;
20'b00001100110000010001 : ColourData = 12'h000;
20'b00001101000000010001 : ColourData = 12'h000;
20'b00001101010000010001 : ColourData = 12'h000;
20'b00001101100000010001 : ColourData = 12'h000;
20'b00001101110000010001 : ColourData = 12'h777;
20'b00001110000000010001 : ColourData = 12'hCCC;
20'b00001110010000010001 : ColourData = 12'hBBB;
20'b00001110100000010001 : ColourData = 12'hBBB;
20'b00001110110000010001 : ColourData = 12'hBBB;
20'b00000000000000010010 : ColourData = 12'h333;
20'b00000000010000010010 : ColourData = 12'h333;
20'b00000000100000010010 : ColourData = 12'h333;
20'b00000000110000010010 : ColourData = 12'h333;
20'b00000001000000010010 : ColourData = 12'h333;
20'b00000001010000010010 : ColourData = 12'h444;
20'b00000001100000010010 : ColourData = 12'h444;
20'b00000001110000010010 : ColourData = 12'h444;
20'b00000010000000010010 : ColourData = 12'h444;
20'b00000010010000010010 : ColourData = 12'h444;
20'b00000010100000010010 : ColourData = 12'h444;
20'b00000010110000010010 : ColourData = 12'h444;
20'b00000011000000010010 : ColourData = 12'h444;
20'b00000011010000010010 : ColourData = 12'h443;
20'b00000011100000010010 : ColourData = 12'h360;
20'b00000011110000010010 : ColourData = 12'h360;
20'b00000100000000010010 : ColourData = 12'h360;
20'b00000100010000010010 : ColourData = 12'h360;
20'b00000100100000010010 : ColourData = 12'h360;
20'b00000100110000010010 : ColourData = 12'h360;
20'b00000101000000010010 : ColourData = 12'h360;
20'b00000101010000010010 : ColourData = 12'h360;
20'b00000101100000010010 : ColourData = 12'h360;
20'b00000101110000010010 : ColourData = 12'h360;
20'b00000110000000010010 : ColourData = 12'h360;
20'b00000110010000010010 : ColourData = 12'h360;
20'b00000110100000010010 : ColourData = 12'h360;
20'b00000110110000010010 : ColourData = 12'h240;
20'b00000111000000010010 : ColourData = 12'h000;
20'b00000111010000010010 : ColourData = 12'h000;
20'b00000111100000010010 : ColourData = 12'h000;
20'b00000111110000010010 : ColourData = 12'h000;
20'b00001000000000010010 : ColourData = 12'h240;
20'b00001000010000010010 : ColourData = 12'h360;
20'b00001000100000010010 : ColourData = 12'h360;
20'b00001000110000010010 : ColourData = 12'h360;
20'b00001001000000010010 : ColourData = 12'h360;
20'b00001001010000010010 : ColourData = 12'h360;
20'b00001001100000010010 : ColourData = 12'h360;
20'b00001001110000010010 : ColourData = 12'h360;
20'b00001010000000010010 : ColourData = 12'h360;
20'b00001010010000010010 : ColourData = 12'h360;
20'b00001010100000010010 : ColourData = 12'h360;
20'b00001010110000010010 : ColourData = 12'h360;
20'b00001011000000010010 : ColourData = 12'h360;
20'b00001011010000010010 : ColourData = 12'h360;
20'b00001011100000010010 : ColourData = 12'h443;
20'b00001011110000010010 : ColourData = 12'h444;
20'b00001100000000010010 : ColourData = 12'h444;
20'b00001100010000010010 : ColourData = 12'h444;
20'b00001100100000010010 : ColourData = 12'h444;
20'b00001100110000010010 : ColourData = 12'h444;
20'b00001101000000010010 : ColourData = 12'h444;
20'b00001101010000010010 : ColourData = 12'h444;
20'b00001101100000010010 : ColourData = 12'h444;
20'b00001101110000010010 : ColourData = 12'h333;
20'b00001110000000010010 : ColourData = 12'h333;
20'b00001110010000010010 : ColourData = 12'h333;
20'b00001110100000010010 : ColourData = 12'h333;
20'b00001110110000010010 : ColourData = 12'h333;
20'b00000000000000010011 : ColourData = 12'h111;
20'b00000000010000010011 : ColourData = 12'h111;
20'b00000000100000010011 : ColourData = 12'h111;
20'b00000000110000010011 : ColourData = 12'h111;
20'b00000001000000010011 : ColourData = 12'h111;
20'b00000001010000010011 : ColourData = 12'h111;
20'b00000001100000010011 : ColourData = 12'h111;
20'b00000001110000010011 : ColourData = 12'h111;
20'b00000010000000010011 : ColourData = 12'h111;
20'b00000010010000010011 : ColourData = 12'h111;
20'b00000010100000010011 : ColourData = 12'h111;
20'b00000010110000010011 : ColourData = 12'h111;
20'b00000011000000010011 : ColourData = 12'h111;
20'b00000011010000010011 : ColourData = 12'h121;
20'b00000011100000010011 : ColourData = 12'h360;
20'b00000011110000010011 : ColourData = 12'h360;
20'b00000100000000010011 : ColourData = 12'h360;
20'b00000100010000010011 : ColourData = 12'h360;
20'b00000100100000010011 : ColourData = 12'h360;
20'b00000100110000010011 : ColourData = 12'h360;
20'b00000101000000010011 : ColourData = 12'h360;
20'b00000101010000010011 : ColourData = 12'h481;
20'b00000101100000010011 : ColourData = 12'h481;
20'b00000101110000010011 : ColourData = 12'h481;
20'b00000110000000010011 : ColourData = 12'h481;
20'b00000110010000010011 : ColourData = 12'h481;
20'b00000110100000010011 : ColourData = 12'h591;
20'b00000110110000010011 : ColourData = 12'h350;
20'b00000111000000010011 : ColourData = 12'h000;
20'b00000111010000010011 : ColourData = 12'h000;
20'b00000111100000010011 : ColourData = 12'h000;
20'b00000111110000010011 : ColourData = 12'h000;
20'b00001000000000010011 : ColourData = 12'h350;
20'b00001000010000010011 : ColourData = 12'h591;
20'b00001000100000010011 : ColourData = 12'h481;
20'b00001000110000010011 : ColourData = 12'h481;
20'b00001001000000010011 : ColourData = 12'h481;
20'b00001001010000010011 : ColourData = 12'h360;
20'b00001001100000010011 : ColourData = 12'h360;
20'b00001001110000010011 : ColourData = 12'h360;
20'b00001010000000010011 : ColourData = 12'h360;
20'b00001010010000010011 : ColourData = 12'h360;
20'b00001010100000010011 : ColourData = 12'h360;
20'b00001010110000010011 : ColourData = 12'h360;
20'b00001011000000010011 : ColourData = 12'h360;
20'b00001011010000010011 : ColourData = 12'h360;
20'b00001011100000010011 : ColourData = 12'h121;
20'b00001011110000010011 : ColourData = 12'h111;
20'b00001100000000010011 : ColourData = 12'h111;
20'b00001100010000010011 : ColourData = 12'h111;
20'b00001100100000010011 : ColourData = 12'h111;
20'b00001100110000010011 : ColourData = 12'h111;
20'b00001101000000010011 : ColourData = 12'h111;
20'b00001101010000010011 : ColourData = 12'h111;
20'b00001101100000010011 : ColourData = 12'h111;
20'b00001101110000010011 : ColourData = 12'h111;
20'b00001110000000010011 : ColourData = 12'h111;
20'b00001110010000010011 : ColourData = 12'h111;
20'b00001110100000010011 : ColourData = 12'h111;
20'b00001110110000010011 : ColourData = 12'h111;
20'b00000000000000010100 : ColourData = 12'h000;
20'b00000000010000010100 : ColourData = 12'h000;
20'b00000000100000010100 : ColourData = 12'h000;
20'b00000000110000010100 : ColourData = 12'h000;
20'b00000001000000010100 : ColourData = 12'h000;
20'b00000001010000010100 : ColourData = 12'h000;
20'b00000001100000010100 : ColourData = 12'h000;
20'b00000001110000010100 : ColourData = 12'h000;
20'b00000010000000010100 : ColourData = 12'h000;
20'b00000010010000010100 : ColourData = 12'h000;
20'b00000010100000010100 : ColourData = 12'h000;
20'b00000010110000010100 : ColourData = 12'h000;
20'b00000011000000010100 : ColourData = 12'h000;
20'b00000011010000010100 : ColourData = 12'h000;
20'b00000011100000010100 : ColourData = 12'h360;
20'b00000011110000010100 : ColourData = 12'h360;
20'b00000100000000010100 : ColourData = 12'h360;
20'b00000100010000010100 : ColourData = 12'h360;
20'b00000100100000010100 : ColourData = 12'h360;
20'b00000100110000010100 : ColourData = 12'h360;
20'b00000101000000010100 : ColourData = 12'h471;
20'b00000101010000010100 : ColourData = 12'h6A1;
20'b00000101100000010100 : ColourData = 12'h5A1;
20'b00000101110000010100 : ColourData = 12'h5A1;
20'b00000110000000010100 : ColourData = 12'h5A1;
20'b00000110010000010100 : ColourData = 12'h5A1;
20'b00000110100000010100 : ColourData = 12'h6A1;
20'b00000110110000010100 : ColourData = 12'h470;
20'b00000111000000010100 : ColourData = 12'h000;
20'b00000111010000010100 : ColourData = 12'h000;
20'b00000111100000010100 : ColourData = 12'h000;
20'b00000111110000010100 : ColourData = 12'h000;
20'b00001000000000010100 : ColourData = 12'h470;
20'b00001000010000010100 : ColourData = 12'h6A1;
20'b00001000100000010100 : ColourData = 12'h5A1;
20'b00001000110000010100 : ColourData = 12'h5A1;
20'b00001001000000010100 : ColourData = 12'h591;
20'b00001001010000010100 : ColourData = 12'h360;
20'b00001001100000010100 : ColourData = 12'h360;
20'b00001001110000010100 : ColourData = 12'h360;
20'b00001010000000010100 : ColourData = 12'h360;
20'b00001010010000010100 : ColourData = 12'h360;
20'b00001010100000010100 : ColourData = 12'h360;
20'b00001010110000010100 : ColourData = 12'h360;
20'b00001011000000010100 : ColourData = 12'h360;
20'b00001011010000010100 : ColourData = 12'h360;
20'b00001011100000010100 : ColourData = 12'h000;
20'b00001011110000010100 : ColourData = 12'h000;
20'b00001100000000010100 : ColourData = 12'h000;
20'b00001100010000010100 : ColourData = 12'h000;
20'b00001100100000010100 : ColourData = 12'h000;
20'b00001100110000010100 : ColourData = 12'h000;
20'b00001101000000010100 : ColourData = 12'h000;
20'b00001101010000010100 : ColourData = 12'h000;
20'b00001101100000010100 : ColourData = 12'h000;
20'b00001101110000010100 : ColourData = 12'h000;
20'b00001110000000010100 : ColourData = 12'h000;
20'b00001110010000010100 : ColourData = 12'h000;
20'b00001110100000010100 : ColourData = 12'h000;
20'b00001110110000010100 : ColourData = 12'h000;
20'b00000000000000010101 : ColourData = 12'h333;
20'b00000000010000010101 : ColourData = 12'h333;
20'b00000000100000010101 : ColourData = 12'h333;
20'b00000000110000010101 : ColourData = 12'h333;
20'b00000001000000010101 : ColourData = 12'h333;
20'b00000001010000010101 : ColourData = 12'h333;
20'b00000001100000010101 : ColourData = 12'h333;
20'b00000001110000010101 : ColourData = 12'h333;
20'b00000010000000010101 : ColourData = 12'h333;
20'b00000010010000010101 : ColourData = 12'h333;
20'b00000010100000010101 : ColourData = 12'h333;
20'b00000010110000010101 : ColourData = 12'h333;
20'b00000011000000010101 : ColourData = 12'h333;
20'b00000011010000010101 : ColourData = 12'h332;
20'b00000011100000010101 : ColourData = 12'h360;
20'b00000011110000010101 : ColourData = 12'h360;
20'b00000100000000010101 : ColourData = 12'h360;
20'b00000100010000010101 : ColourData = 12'h360;
20'b00000100100000010101 : ColourData = 12'h360;
20'b00000100110000010101 : ColourData = 12'h360;
20'b00000101000000010101 : ColourData = 12'h470;
20'b00000101010000010101 : ColourData = 12'h5A1;
20'b00000101100000010101 : ColourData = 12'h5A1;
20'b00000101110000010101 : ColourData = 12'h5A1;
20'b00000110000000010101 : ColourData = 12'h5A1;
20'b00000110010000010101 : ColourData = 12'h5A1;
20'b00000110100000010101 : ColourData = 12'h6A1;
20'b00000110110000010101 : ColourData = 12'h360;
20'b00000111000000010101 : ColourData = 12'h000;
20'b00000111010000010101 : ColourData = 12'h000;
20'b00000111100000010101 : ColourData = 12'h000;
20'b00000111110000010101 : ColourData = 12'h000;
20'b00001000000000010101 : ColourData = 12'h360;
20'b00001000010000010101 : ColourData = 12'h6A1;
20'b00001000100000010101 : ColourData = 12'h5A1;
20'b00001000110000010101 : ColourData = 12'h5A1;
20'b00001001000000010101 : ColourData = 12'h591;
20'b00001001010000010101 : ColourData = 12'h360;
20'b00001001100000010101 : ColourData = 12'h360;
20'b00001001110000010101 : ColourData = 12'h360;
20'b00001010000000010101 : ColourData = 12'h360;
20'b00001010010000010101 : ColourData = 12'h360;
20'b00001010100000010101 : ColourData = 12'h360;
20'b00001010110000010101 : ColourData = 12'h360;
20'b00001011000000010101 : ColourData = 12'h360;
20'b00001011010000010101 : ColourData = 12'h360;
20'b00001011100000010101 : ColourData = 12'h332;
20'b00001011110000010101 : ColourData = 12'h333;
20'b00001100000000010101 : ColourData = 12'h333;
20'b00001100010000010101 : ColourData = 12'h333;
20'b00001100100000010101 : ColourData = 12'h333;
20'b00001100110000010101 : ColourData = 12'h333;
20'b00001101000000010101 : ColourData = 12'h333;
20'b00001101010000010101 : ColourData = 12'h333;
20'b00001101100000010101 : ColourData = 12'h333;
20'b00001101110000010101 : ColourData = 12'h333;
20'b00001110000000010101 : ColourData = 12'h333;
20'b00001110010000010101 : ColourData = 12'h333;
20'b00001110100000010101 : ColourData = 12'h333;
20'b00001110110000010101 : ColourData = 12'h333;
20'b00000000000000010110 : ColourData = 12'h333;
20'b00000000010000010110 : ColourData = 12'h333;
20'b00000000100000010110 : ColourData = 12'h333;
20'b00000000110000010110 : ColourData = 12'h333;
20'b00000001000000010110 : ColourData = 12'h333;
20'b00000001010000010110 : ColourData = 12'h333;
20'b00000001100000010110 : ColourData = 12'h333;
20'b00000001110000010110 : ColourData = 12'h443;
20'b00000010000000010110 : ColourData = 12'h443;
20'b00000010010000010110 : ColourData = 12'h443;
20'b00000010100000010110 : ColourData = 12'h443;
20'b00000010110000010110 : ColourData = 12'h443;
20'b00000011000000010110 : ColourData = 12'h444;
20'b00000011010000010110 : ColourData = 12'h343;
20'b00000011100000010110 : ColourData = 12'h360;
20'b00000011110000010110 : ColourData = 12'h360;
20'b00000100000000010110 : ColourData = 12'h360;
20'b00000100010000010110 : ColourData = 12'h360;
20'b00000100100000010110 : ColourData = 12'h360;
20'b00000100110000010110 : ColourData = 12'h360;
20'b00000101000000010110 : ColourData = 12'h471;
20'b00000101010000010110 : ColourData = 12'h5A1;
20'b00000101100000010110 : ColourData = 12'h5A1;
20'b00000101110000010110 : ColourData = 12'h5A1;
20'b00000110000000010110 : ColourData = 12'h5A1;
20'b00000110010000010110 : ColourData = 12'h5A1;
20'b00000110100000010110 : ColourData = 12'h6A1;
20'b00000110110000010110 : ColourData = 12'h360;
20'b00000111000000010110 : ColourData = 12'h000;
20'b00000111010000010110 : ColourData = 12'h000;
20'b00000111100000010110 : ColourData = 12'h000;
20'b00000111110000010110 : ColourData = 12'h000;
20'b00001000000000010110 : ColourData = 12'h360;
20'b00001000010000010110 : ColourData = 12'h6A1;
20'b00001000100000010110 : ColourData = 12'h5A1;
20'b00001000110000010110 : ColourData = 12'h5A1;
20'b00001001000000010110 : ColourData = 12'h591;
20'b00001001010000010110 : ColourData = 12'h360;
20'b00001001100000010110 : ColourData = 12'h360;
20'b00001001110000010110 : ColourData = 12'h360;
20'b00001010000000010110 : ColourData = 12'h360;
20'b00001010010000010110 : ColourData = 12'h360;
20'b00001010100000010110 : ColourData = 12'h360;
20'b00001010110000010110 : ColourData = 12'h360;
20'b00001011000000010110 : ColourData = 12'h360;
20'b00001011010000010110 : ColourData = 12'h360;
20'b00001011100000010110 : ColourData = 12'h343;
20'b00001011110000010110 : ColourData = 12'h444;
20'b00001100000000010110 : ColourData = 12'h443;
20'b00001100010000010110 : ColourData = 12'h443;
20'b00001100100000010110 : ColourData = 12'h443;
20'b00001100110000010110 : ColourData = 12'h443;
20'b00001101000000010110 : ColourData = 12'h443;
20'b00001101010000010110 : ColourData = 12'h333;
20'b00001101100000010110 : ColourData = 12'h333;
20'b00001101110000010110 : ColourData = 12'h333;
20'b00001110000000010110 : ColourData = 12'h333;
20'b00001110010000010110 : ColourData = 12'h333;
20'b00001110100000010110 : ColourData = 12'h333;
20'b00001110110000010110 : ColourData = 12'h333;
20'b00000000000000010111 : ColourData = 12'h000;
20'b00000000010000010111 : ColourData = 12'h000;
20'b00000000100000010111 : ColourData = 12'h000;
20'b00000000110000010111 : ColourData = 12'h000;
20'b00000001000000010111 : ColourData = 12'h000;
20'b00000001010000010111 : ColourData = 12'h000;
20'b00000001100000010111 : ColourData = 12'h000;
20'b00000001110000010111 : ColourData = 12'h360;
20'b00000010000000010111 : ColourData = 12'h360;
20'b00000010010000010111 : ColourData = 12'h360;
20'b00000010100000010111 : ColourData = 12'h360;
20'b00000010110000010111 : ColourData = 12'h360;
20'b00000011000000010111 : ColourData = 12'h360;
20'b00000011010000010111 : ColourData = 12'h360;
20'b00000011100000010111 : ColourData = 12'h5A1;
20'b00000011110000010111 : ColourData = 12'h5A1;
20'b00000100000000010111 : ColourData = 12'h5A1;
20'b00000100010000010111 : ColourData = 12'h5A1;
20'b00000100100000010111 : ColourData = 12'h5A1;
20'b00000100110000010111 : ColourData = 12'h5A1;
20'b00000101000000010111 : ColourData = 12'h5A1;
20'b00000101010000010111 : ColourData = 12'h5A1;
20'b00000101100000010111 : ColourData = 12'h5A1;
20'b00000101110000010111 : ColourData = 12'h5A1;
20'b00000110000000010111 : ColourData = 12'h5A1;
20'b00000110010000010111 : ColourData = 12'h5A1;
20'b00000110100000010111 : ColourData = 12'h6A1;
20'b00000110110000010111 : ColourData = 12'h360;
20'b00000111000000010111 : ColourData = 12'h000;
20'b00000111010000010111 : ColourData = 12'h000;
20'b00000111100000010111 : ColourData = 12'h000;
20'b00000111110000010111 : ColourData = 12'h000;
20'b00001000000000010111 : ColourData = 12'h360;
20'b00001000010000010111 : ColourData = 12'h6A1;
20'b00001000100000010111 : ColourData = 12'h5A1;
20'b00001000110000010111 : ColourData = 12'h5A1;
20'b00001001000000010111 : ColourData = 12'h5A1;
20'b00001001010000010111 : ColourData = 12'h5A1;
20'b00001001100000010111 : ColourData = 12'h5A1;
20'b00001001110000010111 : ColourData = 12'h5A1;
20'b00001010000000010111 : ColourData = 12'h5A1;
20'b00001010010000010111 : ColourData = 12'h5A1;
20'b00001010100000010111 : ColourData = 12'h5A1;
20'b00001010110000010111 : ColourData = 12'h5A1;
20'b00001011000000010111 : ColourData = 12'h5A1;
20'b00001011010000010111 : ColourData = 12'h5A1;
20'b00001011100000010111 : ColourData = 12'h360;
20'b00001011110000010111 : ColourData = 12'h360;
20'b00001100000000010111 : ColourData = 12'h360;
20'b00001100010000010111 : ColourData = 12'h360;
20'b00001100100000010111 : ColourData = 12'h360;
20'b00001100110000010111 : ColourData = 12'h360;
20'b00001101000000010111 : ColourData = 12'h360;
20'b00001101010000010111 : ColourData = 12'h000;
20'b00001101100000010111 : ColourData = 12'h000;
20'b00001101110000010111 : ColourData = 12'h000;
20'b00001110000000010111 : ColourData = 12'h000;
20'b00001110010000010111 : ColourData = 12'h000;
20'b00001110100000010111 : ColourData = 12'h000;
20'b00001110110000010111 : ColourData = 12'h000;
20'b00000000000000011000 : ColourData = 12'h000;
20'b00000000010000011000 : ColourData = 12'h000;
20'b00000000100000011000 : ColourData = 12'h000;
20'b00000000110000011000 : ColourData = 12'h000;
20'b00000001000000011000 : ColourData = 12'h000;
20'b00000001010000011000 : ColourData = 12'h000;
20'b00000001100000011000 : ColourData = 12'h010;
20'b00000001110000011000 : ColourData = 12'h360;
20'b00000010000000011000 : ColourData = 12'h360;
20'b00000010010000011000 : ColourData = 12'h360;
20'b00000010100000011000 : ColourData = 12'h360;
20'b00000010110000011000 : ColourData = 12'h360;
20'b00000011000000011000 : ColourData = 12'h471;
20'b00000011010000011000 : ColourData = 12'h471;
20'b00000011100000011000 : ColourData = 12'h5A1;
20'b00000011110000011000 : ColourData = 12'h5A1;
20'b00000100000000011000 : ColourData = 12'h5A1;
20'b00000100010000011000 : ColourData = 12'h5A1;
20'b00000100100000011000 : ColourData = 12'h5A1;
20'b00000100110000011000 : ColourData = 12'h5A1;
20'b00000101000000011000 : ColourData = 12'h5A1;
20'b00000101010000011000 : ColourData = 12'h5A1;
20'b00000101100000011000 : ColourData = 12'h5A1;
20'b00000101110000011000 : ColourData = 12'h5A1;
20'b00000110000000011000 : ColourData = 12'h5A1;
20'b00000110010000011000 : ColourData = 12'h5A1;
20'b00000110100000011000 : ColourData = 12'h6A1;
20'b00000110110000011000 : ColourData = 12'h360;
20'b00000111000000011000 : ColourData = 12'h000;
20'b00000111010000011000 : ColourData = 12'h000;
20'b00000111100000011000 : ColourData = 12'h000;
20'b00000111110000011000 : ColourData = 12'h000;
20'b00001000000000011000 : ColourData = 12'h360;
20'b00001000010000011000 : ColourData = 12'h6A1;
20'b00001000100000011000 : ColourData = 12'h5A1;
20'b00001000110000011000 : ColourData = 12'h5A1;
20'b00001001000000011000 : ColourData = 12'h5A1;
20'b00001001010000011000 : ColourData = 12'h5A1;
20'b00001001100000011000 : ColourData = 12'h5A1;
20'b00001001110000011000 : ColourData = 12'h5A1;
20'b00001010000000011000 : ColourData = 12'h5A1;
20'b00001010010000011000 : ColourData = 12'h5A1;
20'b00001010100000011000 : ColourData = 12'h5A1;
20'b00001010110000011000 : ColourData = 12'h5A1;
20'b00001011000000011000 : ColourData = 12'h5A1;
20'b00001011010000011000 : ColourData = 12'h5A1;
20'b00001011100000011000 : ColourData = 12'h471;
20'b00001011110000011000 : ColourData = 12'h471;
20'b00001100000000011000 : ColourData = 12'h360;
20'b00001100010000011000 : ColourData = 12'h360;
20'b00001100100000011000 : ColourData = 12'h360;
20'b00001100110000011000 : ColourData = 12'h360;
20'b00001101000000011000 : ColourData = 12'h360;
20'b00001101010000011000 : ColourData = 12'h010;
20'b00001101100000011000 : ColourData = 12'h000;
20'b00001101110000011000 : ColourData = 12'h000;
20'b00001110000000011000 : ColourData = 12'h000;
20'b00001110010000011000 : ColourData = 12'h000;
20'b00001110100000011000 : ColourData = 12'h000;
20'b00001110110000011000 : ColourData = 12'h000;
20'b00000000000000011001 : ColourData = 12'h444;
20'b00000000010000011001 : ColourData = 12'h444;
20'b00000000100000011001 : ColourData = 12'h444;
20'b00000000110000011001 : ColourData = 12'h444;
20'b00000001000000011001 : ColourData = 12'h444;
20'b00000001010000011001 : ColourData = 12'h444;
20'b00000001100000011001 : ColourData = 12'h444;
20'b00000001110000011001 : ColourData = 12'h360;
20'b00000010000000011001 : ColourData = 12'h360;
20'b00000010010000011001 : ColourData = 12'h360;
20'b00000010100000011001 : ColourData = 12'h350;
20'b00000010110000011001 : ColourData = 12'h481;
20'b00000011000000011001 : ColourData = 12'h6A1;
20'b00000011010000011001 : ColourData = 12'h5A1;
20'b00000011100000011001 : ColourData = 12'h5A1;
20'b00000011110000011001 : ColourData = 12'h5A1;
20'b00000100000000011001 : ColourData = 12'h5A1;
20'b00000100010000011001 : ColourData = 12'h5A1;
20'b00000100100000011001 : ColourData = 12'h5A1;
20'b00000100110000011001 : ColourData = 12'h5A1;
20'b00000101000000011001 : ColourData = 12'h5A1;
20'b00000101010000011001 : ColourData = 12'h5A1;
20'b00000101100000011001 : ColourData = 12'h5A1;
20'b00000101110000011001 : ColourData = 12'h5A1;
20'b00000110000000011001 : ColourData = 12'h5A1;
20'b00000110010000011001 : ColourData = 12'h5A1;
20'b00000110100000011001 : ColourData = 12'h6A1;
20'b00000110110000011001 : ColourData = 12'h470;
20'b00000111000000011001 : ColourData = 12'h000;
20'b00000111010000011001 : ColourData = 12'h000;
20'b00000111100000011001 : ColourData = 12'h000;
20'b00000111110000011001 : ColourData = 12'h000;
20'b00001000000000011001 : ColourData = 12'h470;
20'b00001000010000011001 : ColourData = 12'h6A1;
20'b00001000100000011001 : ColourData = 12'h5A1;
20'b00001000110000011001 : ColourData = 12'h5A1;
20'b00001001000000011001 : ColourData = 12'h5A1;
20'b00001001010000011001 : ColourData = 12'h5A1;
20'b00001001100000011001 : ColourData = 12'h5A1;
20'b00001001110000011001 : ColourData = 12'h5A1;
20'b00001010000000011001 : ColourData = 12'h5A1;
20'b00001010010000011001 : ColourData = 12'h5A1;
20'b00001010100000011001 : ColourData = 12'h5A1;
20'b00001010110000011001 : ColourData = 12'h5A1;
20'b00001011000000011001 : ColourData = 12'h5A1;
20'b00001011010000011001 : ColourData = 12'h5A1;
20'b00001011100000011001 : ColourData = 12'h5A1;
20'b00001011110000011001 : ColourData = 12'h6A1;
20'b00001100000000011001 : ColourData = 12'h481;
20'b00001100010000011001 : ColourData = 12'h350;
20'b00001100100000011001 : ColourData = 12'h360;
20'b00001100110000011001 : ColourData = 12'h360;
20'b00001101000000011001 : ColourData = 12'h360;
20'b00001101010000011001 : ColourData = 12'h444;
20'b00001101100000011001 : ColourData = 12'h444;
20'b00001101110000011001 : ColourData = 12'h444;
20'b00001110000000011001 : ColourData = 12'h444;
20'b00001110010000011001 : ColourData = 12'h444;
20'b00001110100000011001 : ColourData = 12'h444;
20'b00001110110000011001 : ColourData = 12'h444;
20'b00000000000000011010 : ColourData = 12'h111;
20'b00000000010000011010 : ColourData = 12'h111;
20'b00000000100000011010 : ColourData = 12'h111;
20'b00000000110000011010 : ColourData = 12'h111;
20'b00000001000000011010 : ColourData = 12'h111;
20'b00000001010000011010 : ColourData = 12'h111;
20'b00000001100000011010 : ColourData = 12'h121;
20'b00000001110000011010 : ColourData = 12'h360;
20'b00000010000000011010 : ColourData = 12'h360;
20'b00000010010000011010 : ColourData = 12'h471;
20'b00000010100000011010 : ColourData = 12'h481;
20'b00000010110000011010 : ColourData = 12'h591;
20'b00000011000000011010 : ColourData = 12'h5A1;
20'b00000011010000011010 : ColourData = 12'h5A1;
20'b00000011100000011010 : ColourData = 12'h5A1;
20'b00000011110000011010 : ColourData = 12'h5A1;
20'b00000100000000011010 : ColourData = 12'h5A1;
20'b00000100010000011010 : ColourData = 12'h5A1;
20'b00000100100000011010 : ColourData = 12'h581;
20'b00000100110000011010 : ColourData = 12'h471;
20'b00000101000000011010 : ColourData = 12'h481;
20'b00000101010000011010 : ColourData = 12'h481;
20'b00000101100000011010 : ColourData = 12'h481;
20'b00000101110000011010 : ColourData = 12'h481;
20'b00000110000000011010 : ColourData = 12'h481;
20'b00000110010000011010 : ColourData = 12'h481;
20'b00000110100000011010 : ColourData = 12'h481;
20'b00000110110000011010 : ColourData = 12'h350;
20'b00000111000000011010 : ColourData = 12'h000;
20'b00000111010000011010 : ColourData = 12'h000;
20'b00000111100000011010 : ColourData = 12'h000;
20'b00000111110000011010 : ColourData = 12'h000;
20'b00001000000000011010 : ColourData = 12'h350;
20'b00001000010000011010 : ColourData = 12'h481;
20'b00001000100000011010 : ColourData = 12'h481;
20'b00001000110000011010 : ColourData = 12'h481;
20'b00001001000000011010 : ColourData = 12'h481;
20'b00001001010000011010 : ColourData = 12'h481;
20'b00001001100000011010 : ColourData = 12'h481;
20'b00001001110000011010 : ColourData = 12'h481;
20'b00001010000000011010 : ColourData = 12'h471;
20'b00001010010000011010 : ColourData = 12'h581;
20'b00001010100000011010 : ColourData = 12'h5A1;
20'b00001010110000011010 : ColourData = 12'h5A1;
20'b00001011000000011010 : ColourData = 12'h5A1;
20'b00001011010000011010 : ColourData = 12'h5A1;
20'b00001011100000011010 : ColourData = 12'h5A1;
20'b00001011110000011010 : ColourData = 12'h5A1;
20'b00001100000000011010 : ColourData = 12'h591;
20'b00001100010000011010 : ColourData = 12'h481;
20'b00001100100000011010 : ColourData = 12'h471;
20'b00001100110000011010 : ColourData = 12'h360;
20'b00001101000000011010 : ColourData = 12'h360;
20'b00001101010000011010 : ColourData = 12'h121;
20'b00001101100000011010 : ColourData = 12'h111;
20'b00001101110000011010 : ColourData = 12'h111;
20'b00001110000000011010 : ColourData = 12'h111;
20'b00001110010000011010 : ColourData = 12'h111;
20'b00001110100000011010 : ColourData = 12'h111;
20'b00001110110000011010 : ColourData = 12'h111;
20'b00000000000000011011 : ColourData = 12'h000;
20'b00000000010000011011 : ColourData = 12'h000;
20'b00000000100000011011 : ColourData = 12'h000;
20'b00000000110000011011 : ColourData = 12'h000;
20'b00000001000000011011 : ColourData = 12'h000;
20'b00000001010000011011 : ColourData = 12'h000;
20'b00000001100000011011 : ColourData = 12'h000;
20'b00000001110000011011 : ColourData = 12'h360;
20'b00000010000000011011 : ColourData = 12'h360;
20'b00000010010000011011 : ColourData = 12'h591;
20'b00000010100000011011 : ColourData = 12'h6A1;
20'b00000010110000011011 : ColourData = 12'h5A1;
20'b00000011000000011011 : ColourData = 12'h5A1;
20'b00000011010000011011 : ColourData = 12'h5A1;
20'b00000011100000011011 : ColourData = 12'h5A1;
20'b00000011110000011011 : ColourData = 12'h5A1;
20'b00000100000000011011 : ColourData = 12'h5A1;
20'b00000100010000011011 : ColourData = 12'h6A1;
20'b00000100100000011011 : ColourData = 12'h481;
20'b00000100110000011011 : ColourData = 12'h350;
20'b00000101000000011011 : ColourData = 12'h360;
20'b00000101010000011011 : ColourData = 12'h360;
20'b00000101100000011011 : ColourData = 12'h360;
20'b00000101110000011011 : ColourData = 12'h360;
20'b00000110000000011011 : ColourData = 12'h360;
20'b00000110010000011011 : ColourData = 12'h360;
20'b00000110100000011011 : ColourData = 12'h360;
20'b00000110110000011011 : ColourData = 12'h240;
20'b00000111000000011011 : ColourData = 12'h000;
20'b00000111010000011011 : ColourData = 12'h000;
20'b00000111100000011011 : ColourData = 12'h000;
20'b00000111110000011011 : ColourData = 12'h000;
20'b00001000000000011011 : ColourData = 12'h240;
20'b00001000010000011011 : ColourData = 12'h360;
20'b00001000100000011011 : ColourData = 12'h360;
20'b00001000110000011011 : ColourData = 12'h360;
20'b00001001000000011011 : ColourData = 12'h360;
20'b00001001010000011011 : ColourData = 12'h360;
20'b00001001100000011011 : ColourData = 12'h360;
20'b00001001110000011011 : ColourData = 12'h360;
20'b00001010000000011011 : ColourData = 12'h350;
20'b00001010010000011011 : ColourData = 12'h481;
20'b00001010100000011011 : ColourData = 12'h6A1;
20'b00001010110000011011 : ColourData = 12'h5A1;
20'b00001011000000011011 : ColourData = 12'h5A1;
20'b00001011010000011011 : ColourData = 12'h5A1;
20'b00001011100000011011 : ColourData = 12'h5A1;
20'b00001011110000011011 : ColourData = 12'h5A1;
20'b00001100000000011011 : ColourData = 12'h5A1;
20'b00001100010000011011 : ColourData = 12'h6A1;
20'b00001100100000011011 : ColourData = 12'h591;
20'b00001100110000011011 : ColourData = 12'h360;
20'b00001101000000011011 : ColourData = 12'h360;
20'b00001101010000011011 : ColourData = 12'h000;
20'b00001101100000011011 : ColourData = 12'h000;
20'b00001101110000011011 : ColourData = 12'h000;
20'b00001110000000011011 : ColourData = 12'h000;
20'b00001110010000011011 : ColourData = 12'h000;
20'b00001110100000011011 : ColourData = 12'h000;
20'b00001110110000011011 : ColourData = 12'h000;
20'b00000000000000011100 : ColourData = 12'h333;
20'b00000000010000011100 : ColourData = 12'h333;
20'b00000000100000011100 : ColourData = 12'h333;
20'b00000000110000011100 : ColourData = 12'h333;
20'b00000001000000011100 : ColourData = 12'h333;
20'b00000001010000011100 : ColourData = 12'h333;
20'b00000001100000011100 : ColourData = 12'h332;
20'b00000001110000011100 : ColourData = 12'h360;
20'b00000010000000011100 : ColourData = 12'h360;
20'b00000010010000011100 : ColourData = 12'h591;
20'b00000010100000011100 : ColourData = 12'h5A1;
20'b00000010110000011100 : ColourData = 12'h5A1;
20'b00000011000000011100 : ColourData = 12'h5A1;
20'b00000011010000011100 : ColourData = 12'h5A1;
20'b00000011100000011100 : ColourData = 12'h5A1;
20'b00000011110000011100 : ColourData = 12'h5A1;
20'b00000100000000011100 : ColourData = 12'h471;
20'b00000100010000011100 : ColourData = 12'h370;
20'b00000100100000011100 : ColourData = 12'h360;
20'b00000100110000011100 : ColourData = 12'h360;
20'b00000101000000011100 : ColourData = 12'h360;
20'b00000101010000011100 : ColourData = 12'h360;
20'b00000101100000011100 : ColourData = 12'h360;
20'b00000101110000011100 : ColourData = 12'h360;
20'b00000110000000011100 : ColourData = 12'h360;
20'b00000110010000011100 : ColourData = 12'h360;
20'b00000110100000011100 : ColourData = 12'h360;
20'b00000110110000011100 : ColourData = 12'h240;
20'b00000111000000011100 : ColourData = 12'h000;
20'b00000111010000011100 : ColourData = 12'h000;
20'b00000111100000011100 : ColourData = 12'h000;
20'b00000111110000011100 : ColourData = 12'h000;
20'b00001000000000011100 : ColourData = 12'h240;
20'b00001000010000011100 : ColourData = 12'h360;
20'b00001000100000011100 : ColourData = 12'h360;
20'b00001000110000011100 : ColourData = 12'h360;
20'b00001001000000011100 : ColourData = 12'h360;
20'b00001001010000011100 : ColourData = 12'h360;
20'b00001001100000011100 : ColourData = 12'h360;
20'b00001001110000011100 : ColourData = 12'h360;
20'b00001010000000011100 : ColourData = 12'h360;
20'b00001010010000011100 : ColourData = 12'h360;
20'b00001010100000011100 : ColourData = 12'h370;
20'b00001010110000011100 : ColourData = 12'h471;
20'b00001011000000011100 : ColourData = 12'h5A1;
20'b00001011010000011100 : ColourData = 12'h5A1;
20'b00001011100000011100 : ColourData = 12'h5A1;
20'b00001011110000011100 : ColourData = 12'h5A1;
20'b00001100000000011100 : ColourData = 12'h5A1;
20'b00001100010000011100 : ColourData = 12'h5A1;
20'b00001100100000011100 : ColourData = 12'h591;
20'b00001100110000011100 : ColourData = 12'h360;
20'b00001101000000011100 : ColourData = 12'h360;
20'b00001101010000011100 : ColourData = 12'h332;
20'b00001101100000011100 : ColourData = 12'h333;
20'b00001101110000011100 : ColourData = 12'h333;
20'b00001110000000011100 : ColourData = 12'h333;
20'b00001110010000011100 : ColourData = 12'h333;
20'b00001110100000011100 : ColourData = 12'h333;
20'b00001110110000011100 : ColourData = 12'h333;
20'b00000000000000011101 : ColourData = 12'h333;
20'b00000000010000011101 : ColourData = 12'h333;
20'b00000000100000011101 : ColourData = 12'h333;
20'b00000000110000011101 : ColourData = 12'h333;
20'b00000001000000011101 : ColourData = 12'h333;
20'b00000001010000011101 : ColourData = 12'h334;
20'b00000001100000011101 : ColourData = 12'h343;
20'b00000001110000011101 : ColourData = 12'h360;
20'b00000010000000011101 : ColourData = 12'h360;
20'b00000010010000011101 : ColourData = 12'h591;
20'b00000010100000011101 : ColourData = 12'h5A1;
20'b00000010110000011101 : ColourData = 12'h5A1;
20'b00000011000000011101 : ColourData = 12'h5A1;
20'b00000011010000011101 : ColourData = 12'h5A1;
20'b00000011100000011101 : ColourData = 12'h591;
20'b00000011110000011101 : ColourData = 12'h5A1;
20'b00000100000000011101 : ColourData = 12'h360;
20'b00000100010000011101 : ColourData = 12'h360;
20'b00000100100000011101 : ColourData = 12'h360;
20'b00000100110000011101 : ColourData = 12'h360;
20'b00000101000000011101 : ColourData = 12'h360;
20'b00000101010000011101 : ColourData = 12'h360;
20'b00000101100000011101 : ColourData = 12'h360;
20'b00000101110000011101 : ColourData = 12'h360;
20'b00000110000000011101 : ColourData = 12'h360;
20'b00000110010000011101 : ColourData = 12'h360;
20'b00000110100000011101 : ColourData = 12'h360;
20'b00000110110000011101 : ColourData = 12'h240;
20'b00000111000000011101 : ColourData = 12'h000;
20'b00000111010000011101 : ColourData = 12'h000;
20'b00000111100000011101 : ColourData = 12'h000;
20'b00000111110000011101 : ColourData = 12'h000;
20'b00001000000000011101 : ColourData = 12'h240;
20'b00001000010000011101 : ColourData = 12'h360;
20'b00001000100000011101 : ColourData = 12'h360;
20'b00001000110000011101 : ColourData = 12'h360;
20'b00001001000000011101 : ColourData = 12'h360;
20'b00001001010000011101 : ColourData = 12'h360;
20'b00001001100000011101 : ColourData = 12'h360;
20'b00001001110000011101 : ColourData = 12'h360;
20'b00001010000000011101 : ColourData = 12'h360;
20'b00001010010000011101 : ColourData = 12'h360;
20'b00001010100000011101 : ColourData = 12'h360;
20'b00001010110000011101 : ColourData = 12'h360;
20'b00001011000000011101 : ColourData = 12'h5A1;
20'b00001011010000011101 : ColourData = 12'h591;
20'b00001011100000011101 : ColourData = 12'h5A1;
20'b00001011110000011101 : ColourData = 12'h5A1;
20'b00001100000000011101 : ColourData = 12'h5A1;
20'b00001100010000011101 : ColourData = 12'h5A1;
20'b00001100100000011101 : ColourData = 12'h591;
20'b00001100110000011101 : ColourData = 12'h360;
20'b00001101000000011101 : ColourData = 12'h360;
20'b00001101010000011101 : ColourData = 12'h343;
20'b00001101100000011101 : ColourData = 12'h334;
20'b00001101110000011101 : ColourData = 12'h333;
20'b00001110000000011101 : ColourData = 12'h333;
20'b00001110010000011101 : ColourData = 12'h333;
20'b00001110100000011101 : ColourData = 12'h333;
20'b00001110110000011101 : ColourData = 12'h333;
20'b00000000000000011110 : ColourData = 12'h000;
20'b00000000010000011110 : ColourData = 12'h000;
20'b00000000100000011110 : ColourData = 12'h000;
20'b00000000110000011110 : ColourData = 12'h000;
20'b00000001000000011110 : ColourData = 12'h000;
20'b00000001010000011110 : ColourData = 12'h000;
20'b00000001100000011110 : ColourData = 12'h000;
20'b00000001110000011110 : ColourData = 12'h360;
20'b00000010000000011110 : ColourData = 12'h360;
20'b00000010010000011110 : ColourData = 12'h591;
20'b00000010100000011110 : ColourData = 12'h5A1;
20'b00000010110000011110 : ColourData = 12'h5A1;
20'b00000011000000011110 : ColourData = 12'h5A1;
20'b00000011010000011110 : ColourData = 12'h591;
20'b00000011100000011110 : ColourData = 12'h360;
20'b00000011110000011110 : ColourData = 12'h360;
20'b00000100000000011110 : ColourData = 12'h360;
20'b00000100010000011110 : ColourData = 12'h360;
20'b00000100100000011110 : ColourData = 12'h481;
20'b00000100110000011110 : ColourData = 12'h5A1;
20'b00000101000000011110 : ColourData = 12'h591;
20'b00000101010000011110 : ColourData = 12'h591;
20'b00000101100000011110 : ColourData = 12'h591;
20'b00000101110000011110 : ColourData = 12'h591;
20'b00000110000000011110 : ColourData = 12'h591;
20'b00000110010000011110 : ColourData = 12'h591;
20'b00000110100000011110 : ColourData = 12'h6A1;
20'b00000110110000011110 : ColourData = 12'h360;
20'b00000111000000011110 : ColourData = 12'h000;
20'b00000111010000011110 : ColourData = 12'h000;
20'b00000111100000011110 : ColourData = 12'h000;
20'b00000111110000011110 : ColourData = 12'h000;
20'b00001000000000011110 : ColourData = 12'h360;
20'b00001000010000011110 : ColourData = 12'h6A1;
20'b00001000100000011110 : ColourData = 12'h591;
20'b00001000110000011110 : ColourData = 12'h591;
20'b00001001000000011110 : ColourData = 12'h591;
20'b00001001010000011110 : ColourData = 12'h591;
20'b00001001100000011110 : ColourData = 12'h591;
20'b00001001110000011110 : ColourData = 12'h591;
20'b00001010000000011110 : ColourData = 12'h5A1;
20'b00001010010000011110 : ColourData = 12'h481;
20'b00001010100000011110 : ColourData = 12'h360;
20'b00001010110000011110 : ColourData = 12'h360;
20'b00001011000000011110 : ColourData = 12'h360;
20'b00001011010000011110 : ColourData = 12'h360;
20'b00001011100000011110 : ColourData = 12'h591;
20'b00001011110000011110 : ColourData = 12'h5A1;
20'b00001100000000011110 : ColourData = 12'h5A1;
20'b00001100010000011110 : ColourData = 12'h5A1;
20'b00001100100000011110 : ColourData = 12'h591;
20'b00001100110000011110 : ColourData = 12'h360;
20'b00001101000000011110 : ColourData = 12'h360;
20'b00001101010000011110 : ColourData = 12'h000;
20'b00001101100000011110 : ColourData = 12'h000;
20'b00001101110000011110 : ColourData = 12'h000;
20'b00001110000000011110 : ColourData = 12'h000;
20'b00001110010000011110 : ColourData = 12'h000;
20'b00001110100000011110 : ColourData = 12'h000;
20'b00001110110000011110 : ColourData = 12'h000;
20'b00000000000000011111 : ColourData = 12'h000;
20'b00000000010000011111 : ColourData = 12'h000;
20'b00000000100000011111 : ColourData = 12'h000;
20'b00000000110000011111 : ColourData = 12'h000;
20'b00000001000000011111 : ColourData = 12'h000;
20'b00000001010000011111 : ColourData = 12'h000;
20'b00000001100000011111 : ColourData = 12'h000;
20'b00000001110000011111 : ColourData = 12'h360;
20'b00000010000000011111 : ColourData = 12'h360;
20'b00000010010000011111 : ColourData = 12'h591;
20'b00000010100000011111 : ColourData = 12'h5A1;
20'b00000010110000011111 : ColourData = 12'h5A1;
20'b00000011000000011111 : ColourData = 12'h5A1;
20'b00000011010000011111 : ColourData = 12'h591;
20'b00000011100000011111 : ColourData = 12'h360;
20'b00000011110000011111 : ColourData = 12'h360;
20'b00000100000000011111 : ColourData = 12'h360;
20'b00000100010000011111 : ColourData = 12'h360;
20'b00000100100000011111 : ColourData = 12'h481;
20'b00000100110000011111 : ColourData = 12'h5A1;
20'b00000101000000011111 : ColourData = 12'h5A1;
20'b00000101010000011111 : ColourData = 12'h5A1;
20'b00000101100000011111 : ColourData = 12'h5A1;
20'b00000101110000011111 : ColourData = 12'h5A1;
20'b00000110000000011111 : ColourData = 12'h5A1;
20'b00000110010000011111 : ColourData = 12'h5A1;
20'b00000110100000011111 : ColourData = 12'h6A1;
20'b00000110110000011111 : ColourData = 12'h471;
20'b00000111000000011111 : ColourData = 12'h010;
20'b00000111010000011111 : ColourData = 12'h010;
20'b00000111100000011111 : ColourData = 12'h010;
20'b00000111110000011111 : ColourData = 12'h010;
20'b00001000000000011111 : ColourData = 12'h471;
20'b00001000010000011111 : ColourData = 12'h6A1;
20'b00001000100000011111 : ColourData = 12'h5A1;
20'b00001000110000011111 : ColourData = 12'h5A1;
20'b00001001000000011111 : ColourData = 12'h5A1;
20'b00001001010000011111 : ColourData = 12'h5A1;
20'b00001001100000011111 : ColourData = 12'h5A1;
20'b00001001110000011111 : ColourData = 12'h5A1;
20'b00001010000000011111 : ColourData = 12'h5A1;
20'b00001010010000011111 : ColourData = 12'h481;
20'b00001010100000011111 : ColourData = 12'h360;
20'b00001010110000011111 : ColourData = 12'h360;
20'b00001011000000011111 : ColourData = 12'h360;
20'b00001011010000011111 : ColourData = 12'h360;
20'b00001011100000011111 : ColourData = 12'h591;
20'b00001011110000011111 : ColourData = 12'h5A1;
20'b00001100000000011111 : ColourData = 12'h5A1;
20'b00001100010000011111 : ColourData = 12'h5A1;
20'b00001100100000011111 : ColourData = 12'h591;
20'b00001100110000011111 : ColourData = 12'h360;
20'b00001101000000011111 : ColourData = 12'h360;
20'b00001101010000011111 : ColourData = 12'h000;
20'b00001101100000011111 : ColourData = 12'h000;
20'b00001101110000011111 : ColourData = 12'h000;
20'b00001110000000011111 : ColourData = 12'h000;
20'b00001110010000011111 : ColourData = 12'h000;
20'b00001110100000011111 : ColourData = 12'h000;
20'b00001110110000011111 : ColourData = 12'h000;
20'b00000000000000100000 : ColourData = 12'h444;
20'b00000000010000100000 : ColourData = 12'h444;
20'b00000000100000100000 : ColourData = 12'h444;
20'b00000000110000100000 : ColourData = 12'h444;
20'b00000001000000100000 : ColourData = 12'h444;
20'b00000001010000100000 : ColourData = 12'h444;
20'b00000001100000100000 : ColourData = 12'h444;
20'b00000001110000100000 : ColourData = 12'h360;
20'b00000010000000100000 : ColourData = 12'h360;
20'b00000010010000100000 : ColourData = 12'h591;
20'b00000010100000100000 : ColourData = 12'h5A1;
20'b00000010110000100000 : ColourData = 12'h5A1;
20'b00000011000000100000 : ColourData = 12'h5A1;
20'b00000011010000100000 : ColourData = 12'h591;
20'b00000011100000100000 : ColourData = 12'h360;
20'b00000011110000100000 : ColourData = 12'h360;
20'b00000100000000100000 : ColourData = 12'h360;
20'b00000100010000100000 : ColourData = 12'h360;
20'b00000100100000100000 : ColourData = 12'h481;
20'b00000100110000100000 : ColourData = 12'h5A1;
20'b00000101000000100000 : ColourData = 12'h5A1;
20'b00000101010000100000 : ColourData = 12'h5A1;
20'b00000101100000100000 : ColourData = 12'h5A1;
20'b00000101110000100000 : ColourData = 12'h5A1;
20'b00000110000000100000 : ColourData = 12'h5A1;
20'b00000110010000100000 : ColourData = 12'h5A1;
20'b00000110100000100000 : ColourData = 12'h591;
20'b00000110110000100000 : ColourData = 12'h5A1;
20'b00000111000000100000 : ColourData = 12'h6A1;
20'b00000111010000100000 : ColourData = 12'h6A1;
20'b00000111100000100000 : ColourData = 12'h6A1;
20'b00000111110000100000 : ColourData = 12'h6A1;
20'b00001000000000100000 : ColourData = 12'h5A1;
20'b00001000010000100000 : ColourData = 12'h591;
20'b00001000100000100000 : ColourData = 12'h5A1;
20'b00001000110000100000 : ColourData = 12'h5A1;
20'b00001001000000100000 : ColourData = 12'h5A1;
20'b00001001010000100000 : ColourData = 12'h5A1;
20'b00001001100000100000 : ColourData = 12'h5A1;
20'b00001001110000100000 : ColourData = 12'h5A1;
20'b00001010000000100000 : ColourData = 12'h5A1;
20'b00001010010000100000 : ColourData = 12'h481;
20'b00001010100000100000 : ColourData = 12'h360;
20'b00001010110000100000 : ColourData = 12'h360;
20'b00001011000000100000 : ColourData = 12'h360;
20'b00001011010000100000 : ColourData = 12'h360;
20'b00001011100000100000 : ColourData = 12'h591;
20'b00001011110000100000 : ColourData = 12'h5A1;
20'b00001100000000100000 : ColourData = 12'h5A1;
20'b00001100010000100000 : ColourData = 12'h5A1;
20'b00001100100000100000 : ColourData = 12'h591;
20'b00001100110000100000 : ColourData = 12'h360;
20'b00001101000000100000 : ColourData = 12'h360;
20'b00001101010000100000 : ColourData = 12'h444;
20'b00001101100000100000 : ColourData = 12'h444;
20'b00001101110000100000 : ColourData = 12'h444;
20'b00001110000000100000 : ColourData = 12'h444;
20'b00001110010000100000 : ColourData = 12'h444;
20'b00001110100000100000 : ColourData = 12'h444;
20'b00001110110000100000 : ColourData = 12'h444;
20'b00000000000000100001 : ColourData = 12'h111;
20'b00000000010000100001 : ColourData = 12'h111;
20'b00000000100000100001 : ColourData = 12'h111;
20'b00000000110000100001 : ColourData = 12'h111;
20'b00000001000000100001 : ColourData = 12'h111;
20'b00000001010000100001 : ColourData = 12'h111;
20'b00000001100000100001 : ColourData = 12'h221;
20'b00000001110000100001 : ColourData = 12'h360;
20'b00000010000000100001 : ColourData = 12'h360;
20'b00000010010000100001 : ColourData = 12'h591;
20'b00000010100000100001 : ColourData = 12'h5A1;
20'b00000010110000100001 : ColourData = 12'h5A1;
20'b00000011000000100001 : ColourData = 12'h5A1;
20'b00000011010000100001 : ColourData = 12'h591;
20'b00000011100000100001 : ColourData = 12'h360;
20'b00000011110000100001 : ColourData = 12'h360;
20'b00000100000000100001 : ColourData = 12'h360;
20'b00000100010000100001 : ColourData = 12'h360;
20'b00000100100000100001 : ColourData = 12'h481;
20'b00000100110000100001 : ColourData = 12'h5A1;
20'b00000101000000100001 : ColourData = 12'h5A1;
20'b00000101010000100001 : ColourData = 12'h5A1;
20'b00000101100000100001 : ColourData = 12'h5A1;
20'b00000101110000100001 : ColourData = 12'h5A1;
20'b00000110000000100001 : ColourData = 12'h5A1;
20'b00000110010000100001 : ColourData = 12'h5A1;
20'b00000110100000100001 : ColourData = 12'h5A1;
20'b00000110110000100001 : ColourData = 12'h5A1;
20'b00000111000000100001 : ColourData = 12'h5A1;
20'b00000111010000100001 : ColourData = 12'h5A1;
20'b00000111100000100001 : ColourData = 12'h5A1;
20'b00000111110000100001 : ColourData = 12'h5A1;
20'b00001000000000100001 : ColourData = 12'h5A1;
20'b00001000010000100001 : ColourData = 12'h5A1;
20'b00001000100000100001 : ColourData = 12'h5A1;
20'b00001000110000100001 : ColourData = 12'h5A1;
20'b00001001000000100001 : ColourData = 12'h5A1;
20'b00001001010000100001 : ColourData = 12'h5A1;
20'b00001001100000100001 : ColourData = 12'h5A1;
20'b00001001110000100001 : ColourData = 12'h5A1;
20'b00001010000000100001 : ColourData = 12'h5A1;
20'b00001010010000100001 : ColourData = 12'h481;
20'b00001010100000100001 : ColourData = 12'h360;
20'b00001010110000100001 : ColourData = 12'h360;
20'b00001011000000100001 : ColourData = 12'h360;
20'b00001011010000100001 : ColourData = 12'h360;
20'b00001011100000100001 : ColourData = 12'h591;
20'b00001011110000100001 : ColourData = 12'h5A1;
20'b00001100000000100001 : ColourData = 12'h5A1;
20'b00001100010000100001 : ColourData = 12'h5A1;
20'b00001100100000100001 : ColourData = 12'h591;
20'b00001100110000100001 : ColourData = 12'h360;
20'b00001101000000100001 : ColourData = 12'h360;
20'b00001101010000100001 : ColourData = 12'h221;
20'b00001101100000100001 : ColourData = 12'h111;
20'b00001101110000100001 : ColourData = 12'h111;
20'b00001110000000100001 : ColourData = 12'h111;
20'b00001110010000100001 : ColourData = 12'h111;
20'b00001110100000100001 : ColourData = 12'h111;
20'b00001110110000100001 : ColourData = 12'h111;
20'b00000000000000100010 : ColourData = 12'h000;
20'b00000000010000100010 : ColourData = 12'h000;
20'b00000000100000100010 : ColourData = 12'h000;
20'b00000000110000100010 : ColourData = 12'h000;
20'b00000001000000100010 : ColourData = 12'h000;
20'b00000001010000100010 : ColourData = 12'h000;
20'b00000001100000100010 : ColourData = 12'h000;
20'b00000001110000100010 : ColourData = 12'h360;
20'b00000010000000100010 : ColourData = 12'h360;
20'b00000010010000100010 : ColourData = 12'h591;
20'b00000010100000100010 : ColourData = 12'h5A1;
20'b00000010110000100010 : ColourData = 12'h5A1;
20'b00000011000000100010 : ColourData = 12'h5A1;
20'b00000011010000100010 : ColourData = 12'h591;
20'b00000011100000100010 : ColourData = 12'h360;
20'b00000011110000100010 : ColourData = 12'h360;
20'b00000100000000100010 : ColourData = 12'h360;
20'b00000100010000100010 : ColourData = 12'h360;
20'b00000100100000100010 : ColourData = 12'h481;
20'b00000100110000100010 : ColourData = 12'h5A1;
20'b00000101000000100010 : ColourData = 12'h5A1;
20'b00000101010000100010 : ColourData = 12'h5A1;
20'b00000101100000100010 : ColourData = 12'h5A1;
20'b00000101110000100010 : ColourData = 12'h5A1;
20'b00000110000000100010 : ColourData = 12'h5A1;
20'b00000110010000100010 : ColourData = 12'h5A1;
20'b00000110100000100010 : ColourData = 12'h5A1;
20'b00000110110000100010 : ColourData = 12'h5A1;
20'b00000111000000100010 : ColourData = 12'h5A1;
20'b00000111010000100010 : ColourData = 12'h5A1;
20'b00000111100000100010 : ColourData = 12'h5A1;
20'b00000111110000100010 : ColourData = 12'h5A1;
20'b00001000000000100010 : ColourData = 12'h5A1;
20'b00001000010000100010 : ColourData = 12'h5A1;
20'b00001000100000100010 : ColourData = 12'h5A1;
20'b00001000110000100010 : ColourData = 12'h5A1;
20'b00001001000000100010 : ColourData = 12'h5A1;
20'b00001001010000100010 : ColourData = 12'h5A1;
20'b00001001100000100010 : ColourData = 12'h5A1;
20'b00001001110000100010 : ColourData = 12'h5A1;
20'b00001010000000100010 : ColourData = 12'h5A1;
20'b00001010010000100010 : ColourData = 12'h481;
20'b00001010100000100010 : ColourData = 12'h360;
20'b00001010110000100010 : ColourData = 12'h360;
20'b00001011000000100010 : ColourData = 12'h360;
20'b00001011010000100010 : ColourData = 12'h360;
20'b00001011100000100010 : ColourData = 12'h591;
20'b00001011110000100010 : ColourData = 12'h5A1;
20'b00001100000000100010 : ColourData = 12'h5A1;
20'b00001100010000100010 : ColourData = 12'h5A1;
20'b00001100100000100010 : ColourData = 12'h591;
20'b00001100110000100010 : ColourData = 12'h360;
20'b00001101000000100010 : ColourData = 12'h360;
20'b00001101010000100010 : ColourData = 12'h000;
20'b00001101100000100010 : ColourData = 12'h000;
20'b00001101110000100010 : ColourData = 12'h000;
20'b00001110000000100010 : ColourData = 12'h000;
20'b00001110010000100010 : ColourData = 12'h000;
20'b00001110100000100010 : ColourData = 12'h000;
20'b00001110110000100010 : ColourData = 12'h000;
20'b00000000000000100011 : ColourData = 12'h222;
20'b00000000010000100011 : ColourData = 12'h222;
20'b00000000100000100011 : ColourData = 12'h222;
20'b00000000110000100011 : ColourData = 12'h222;
20'b00000001000000100011 : ColourData = 12'h222;
20'b00000001010000100011 : ColourData = 12'h222;
20'b00000001100000100011 : ColourData = 12'h232;
20'b00000001110000100011 : ColourData = 12'h360;
20'b00000010000000100011 : ColourData = 12'h360;
20'b00000010010000100011 : ColourData = 12'h591;
20'b00000010100000100011 : ColourData = 12'h5A1;
20'b00000010110000100011 : ColourData = 12'h5A1;
20'b00000011000000100011 : ColourData = 12'h5A1;
20'b00000011010000100011 : ColourData = 12'h591;
20'b00000011100000100011 : ColourData = 12'h360;
20'b00000011110000100011 : ColourData = 12'h360;
20'b00000100000000100011 : ColourData = 12'h360;
20'b00000100010000100011 : ColourData = 12'h360;
20'b00000100100000100011 : ColourData = 12'h481;
20'b00000100110000100011 : ColourData = 12'h5A1;
20'b00000101000000100011 : ColourData = 12'h5A1;
20'b00000101010000100011 : ColourData = 12'h5A1;
20'b00000101100000100011 : ColourData = 12'h5A1;
20'b00000101110000100011 : ColourData = 12'h5A1;
20'b00000110000000100011 : ColourData = 12'h5A1;
20'b00000110010000100011 : ColourData = 12'h5A1;
20'b00000110100000100011 : ColourData = 12'h5A1;
20'b00000110110000100011 : ColourData = 12'h5A1;
20'b00000111000000100011 : ColourData = 12'h5A1;
20'b00000111010000100011 : ColourData = 12'h5A1;
20'b00000111100000100011 : ColourData = 12'h5A1;
20'b00000111110000100011 : ColourData = 12'h5A1;
20'b00001000000000100011 : ColourData = 12'h5A1;
20'b00001000010000100011 : ColourData = 12'h5A1;
20'b00001000100000100011 : ColourData = 12'h5A1;
20'b00001000110000100011 : ColourData = 12'h5A1;
20'b00001001000000100011 : ColourData = 12'h5A1;
20'b00001001010000100011 : ColourData = 12'h5A1;
20'b00001001100000100011 : ColourData = 12'h5A1;
20'b00001001110000100011 : ColourData = 12'h5A1;
20'b00001010000000100011 : ColourData = 12'h5A1;
20'b00001010010000100011 : ColourData = 12'h481;
20'b00001010100000100011 : ColourData = 12'h360;
20'b00001010110000100011 : ColourData = 12'h360;
20'b00001011000000100011 : ColourData = 12'h360;
20'b00001011010000100011 : ColourData = 12'h360;
20'b00001011100000100011 : ColourData = 12'h591;
20'b00001011110000100011 : ColourData = 12'h5A1;
20'b00001100000000100011 : ColourData = 12'h5A1;
20'b00001100010000100011 : ColourData = 12'h5A1;
20'b00001100100000100011 : ColourData = 12'h591;
20'b00001100110000100011 : ColourData = 12'h360;
20'b00001101000000100011 : ColourData = 12'h360;
20'b00001101010000100011 : ColourData = 12'h232;
20'b00001101100000100011 : ColourData = 12'h222;
20'b00001101110000100011 : ColourData = 12'h222;
20'b00001110000000100011 : ColourData = 12'h222;
20'b00001110010000100011 : ColourData = 12'h222;
20'b00001110100000100011 : ColourData = 12'h222;
20'b00001110110000100011 : ColourData = 12'h222;
20'b00000000000000100100 : ColourData = 12'h444;
20'b00000000010000100100 : ColourData = 12'h444;
20'b00000000100000100100 : ColourData = 12'h444;
20'b00000000110000100100 : ColourData = 12'h444;
20'b00000001000000100100 : ColourData = 12'h444;
20'b00000001010000100100 : ColourData = 12'h444;
20'b00000001100000100100 : ColourData = 12'h443;
20'b00000001110000100100 : ColourData = 12'h360;
20'b00000010000000100100 : ColourData = 12'h360;
20'b00000010010000100100 : ColourData = 12'h591;
20'b00000010100000100100 : ColourData = 12'h5A1;
20'b00000010110000100100 : ColourData = 12'h5A1;
20'b00000011000000100100 : ColourData = 12'h5A1;
20'b00000011010000100100 : ColourData = 12'h591;
20'b00000011100000100100 : ColourData = 12'h360;
20'b00000011110000100100 : ColourData = 12'h360;
20'b00000100000000100100 : ColourData = 12'h360;
20'b00000100010000100100 : ColourData = 12'h360;
20'b00000100100000100100 : ColourData = 12'h481;
20'b00000100110000100100 : ColourData = 12'h5A1;
20'b00000101000000100100 : ColourData = 12'h5A1;
20'b00000101010000100100 : ColourData = 12'h5A1;
20'b00000101100000100100 : ColourData = 12'h5A1;
20'b00000101110000100100 : ColourData = 12'h5A1;
20'b00000110000000100100 : ColourData = 12'h5A1;
20'b00000110010000100100 : ColourData = 12'h5A1;
20'b00000110100000100100 : ColourData = 12'h5A1;
20'b00000110110000100100 : ColourData = 12'h5A1;
20'b00000111000000100100 : ColourData = 12'h5A1;
20'b00000111010000100100 : ColourData = 12'h5A1;
20'b00000111100000100100 : ColourData = 12'h5A1;
20'b00000111110000100100 : ColourData = 12'h5A1;
20'b00001000000000100100 : ColourData = 12'h5A1;
20'b00001000010000100100 : ColourData = 12'h5A1;
20'b00001000100000100100 : ColourData = 12'h5A1;
20'b00001000110000100100 : ColourData = 12'h5A1;
20'b00001001000000100100 : ColourData = 12'h5A1;
20'b00001001010000100100 : ColourData = 12'h5A1;
20'b00001001100000100100 : ColourData = 12'h5A1;
20'b00001001110000100100 : ColourData = 12'h5A1;
20'b00001010000000100100 : ColourData = 12'h5A1;
20'b00001010010000100100 : ColourData = 12'h481;
20'b00001010100000100100 : ColourData = 12'h360;
20'b00001010110000100100 : ColourData = 12'h360;
20'b00001011000000100100 : ColourData = 12'h360;
20'b00001011010000100100 : ColourData = 12'h360;
20'b00001011100000100100 : ColourData = 12'h591;
20'b00001011110000100100 : ColourData = 12'h5A1;
20'b00001100000000100100 : ColourData = 12'h5A1;
20'b00001100010000100100 : ColourData = 12'h5A1;
20'b00001100100000100100 : ColourData = 12'h591;
20'b00001100110000100100 : ColourData = 12'h360;
20'b00001101000000100100 : ColourData = 12'h360;
20'b00001101010000100100 : ColourData = 12'h443;
20'b00001101100000100100 : ColourData = 12'h444;
20'b00001101110000100100 : ColourData = 12'h444;
20'b00001110000000100100 : ColourData = 12'h444;
20'b00001110010000100100 : ColourData = 12'h444;
20'b00001110100000100100 : ColourData = 12'h444;
20'b00001110110000100100 : ColourData = 12'h444;
20'b00000000000000100101 : ColourData = 12'h000;
20'b00000000010000100101 : ColourData = 12'h000;
20'b00000000100000100101 : ColourData = 12'h000;
20'b00000000110000100101 : ColourData = 12'h000;
20'b00000001000000100101 : ColourData = 12'h000;
20'b00000001010000100101 : ColourData = 12'h000;
20'b00000001100000100101 : ColourData = 12'h000;
20'b00000001110000100101 : ColourData = 12'h360;
20'b00000010000000100101 : ColourData = 12'h360;
20'b00000010010000100101 : ColourData = 12'h591;
20'b00000010100000100101 : ColourData = 12'h5A1;
20'b00000010110000100101 : ColourData = 12'h5A1;
20'b00000011000000100101 : ColourData = 12'h5A1;
20'b00000011010000100101 : ColourData = 12'h591;
20'b00000011100000100101 : ColourData = 12'h360;
20'b00000011110000100101 : ColourData = 12'h360;
20'b00000100000000100101 : ColourData = 12'h360;
20'b00000100010000100101 : ColourData = 12'h360;
20'b00000100100000100101 : ColourData = 12'h481;
20'b00000100110000100101 : ColourData = 12'h5A1;
20'b00000101000000100101 : ColourData = 12'h5A1;
20'b00000101010000100101 : ColourData = 12'h5A1;
20'b00000101100000100101 : ColourData = 12'h5A1;
20'b00000101110000100101 : ColourData = 12'h5A1;
20'b00000110000000100101 : ColourData = 12'h5A1;
20'b00000110010000100101 : ColourData = 12'h5A1;
20'b00000110100000100101 : ColourData = 12'h5A1;
20'b00000110110000100101 : ColourData = 12'h5A1;
20'b00000111000000100101 : ColourData = 12'h5A1;
20'b00000111010000100101 : ColourData = 12'h5A1;
20'b00000111100000100101 : ColourData = 12'h5A1;
20'b00000111110000100101 : ColourData = 12'h5A1;
20'b00001000000000100101 : ColourData = 12'h5A1;
20'b00001000010000100101 : ColourData = 12'h5A1;
20'b00001000100000100101 : ColourData = 12'h5A1;
20'b00001000110000100101 : ColourData = 12'h5A1;
20'b00001001000000100101 : ColourData = 12'h5A1;
20'b00001001010000100101 : ColourData = 12'h5A1;
20'b00001001100000100101 : ColourData = 12'h5A1;
20'b00001001110000100101 : ColourData = 12'h5A1;
20'b00001010000000100101 : ColourData = 12'h5A1;
20'b00001010010000100101 : ColourData = 12'h481;
20'b00001010100000100101 : ColourData = 12'h360;
20'b00001010110000100101 : ColourData = 12'h360;
20'b00001011000000100101 : ColourData = 12'h360;
20'b00001011010000100101 : ColourData = 12'h360;
20'b00001011100000100101 : ColourData = 12'h591;
20'b00001011110000100101 : ColourData = 12'h5A1;
20'b00001100000000100101 : ColourData = 12'h5A1;
20'b00001100010000100101 : ColourData = 12'h5A1;
20'b00001100100000100101 : ColourData = 12'h591;
20'b00001100110000100101 : ColourData = 12'h360;
20'b00001101000000100101 : ColourData = 12'h360;
20'b00001101010000100101 : ColourData = 12'h000;
20'b00001101100000100101 : ColourData = 12'h000;
20'b00001101110000100101 : ColourData = 12'h000;
20'b00001110000000100101 : ColourData = 12'h000;
20'b00001110010000100101 : ColourData = 12'h000;
20'b00001110100000100101 : ColourData = 12'h000;
20'b00001110110000100101 : ColourData = 12'h000;
20'b00000000000000100110 : ColourData = 12'h000;
20'b00000000010000100110 : ColourData = 12'h000;
20'b00000000100000100110 : ColourData = 12'h000;
20'b00000000110000100110 : ColourData = 12'h000;
20'b00000001000000100110 : ColourData = 12'h000;
20'b00000001010000100110 : ColourData = 12'h000;
20'b00000001100000100110 : ColourData = 12'h000;
20'b00000001110000100110 : ColourData = 12'h360;
20'b00000010000000100110 : ColourData = 12'h360;
20'b00000010010000100110 : ColourData = 12'h591;
20'b00000010100000100110 : ColourData = 12'h5A1;
20'b00000010110000100110 : ColourData = 12'h5A1;
20'b00000011000000100110 : ColourData = 12'h5A1;
20'b00000011010000100110 : ColourData = 12'h591;
20'b00000011100000100110 : ColourData = 12'h360;
20'b00000011110000100110 : ColourData = 12'h360;
20'b00000100000000100110 : ColourData = 12'h360;
20'b00000100010000100110 : ColourData = 12'h360;
20'b00000100100000100110 : ColourData = 12'h481;
20'b00000100110000100110 : ColourData = 12'h5A1;
20'b00000101000000100110 : ColourData = 12'h5A1;
20'b00000101010000100110 : ColourData = 12'h5A1;
20'b00000101100000100110 : ColourData = 12'h5A1;
20'b00000101110000100110 : ColourData = 12'h5A1;
20'b00000110000000100110 : ColourData = 12'h5A1;
20'b00000110010000100110 : ColourData = 12'h5A1;
20'b00000110100000100110 : ColourData = 12'h5A1;
20'b00000110110000100110 : ColourData = 12'h5A1;
20'b00000111000000100110 : ColourData = 12'h5A1;
20'b00000111010000100110 : ColourData = 12'h5A1;
20'b00000111100000100110 : ColourData = 12'h5A1;
20'b00000111110000100110 : ColourData = 12'h5A1;
20'b00001000000000100110 : ColourData = 12'h5A1;
20'b00001000010000100110 : ColourData = 12'h5A1;
20'b00001000100000100110 : ColourData = 12'h5A1;
20'b00001000110000100110 : ColourData = 12'h5A1;
20'b00001001000000100110 : ColourData = 12'h5A1;
20'b00001001010000100110 : ColourData = 12'h5A1;
20'b00001001100000100110 : ColourData = 12'h5A1;
20'b00001001110000100110 : ColourData = 12'h5A1;
20'b00001010000000100110 : ColourData = 12'h5A1;
20'b00001010010000100110 : ColourData = 12'h481;
20'b00001010100000100110 : ColourData = 12'h360;
20'b00001010110000100110 : ColourData = 12'h360;
20'b00001011000000100110 : ColourData = 12'h360;
20'b00001011010000100110 : ColourData = 12'h360;
20'b00001011100000100110 : ColourData = 12'h591;
20'b00001011110000100110 : ColourData = 12'h5A1;
20'b00001100000000100110 : ColourData = 12'h5A1;
20'b00001100010000100110 : ColourData = 12'h5A1;
20'b00001100100000100110 : ColourData = 12'h591;
20'b00001100110000100110 : ColourData = 12'h360;
20'b00001101000000100110 : ColourData = 12'h360;
20'b00001101010000100110 : ColourData = 12'h000;
20'b00001101100000100110 : ColourData = 12'h000;
20'b00001101110000100110 : ColourData = 12'h000;
20'b00001110000000100110 : ColourData = 12'h000;
20'b00001110010000100110 : ColourData = 12'h000;
20'b00001110100000100110 : ColourData = 12'h000;
20'b00001110110000100110 : ColourData = 12'h000;
20'b00000000000000100111 : ColourData = 12'h444;
20'b00000000010000100111 : ColourData = 12'h444;
20'b00000000100000100111 : ColourData = 12'h444;
20'b00000000110000100111 : ColourData = 12'h444;
20'b00000001000000100111 : ColourData = 12'h444;
20'b00000001010000100111 : ColourData = 12'h444;
20'b00000001100000100111 : ColourData = 12'h443;
20'b00000001110000100111 : ColourData = 12'h360;
20'b00000010000000100111 : ColourData = 12'h360;
20'b00000010010000100111 : ColourData = 12'h591;
20'b00000010100000100111 : ColourData = 12'h5A1;
20'b00000010110000100111 : ColourData = 12'h5A1;
20'b00000011000000100111 : ColourData = 12'h5A1;
20'b00000011010000100111 : ColourData = 12'h591;
20'b00000011100000100111 : ColourData = 12'h360;
20'b00000011110000100111 : ColourData = 12'h360;
20'b00000100000000100111 : ColourData = 12'h360;
20'b00000100010000100111 : ColourData = 12'h360;
20'b00000100100000100111 : ColourData = 12'h481;
20'b00000100110000100111 : ColourData = 12'h5A1;
20'b00000101000000100111 : ColourData = 12'h5A1;
20'b00000101010000100111 : ColourData = 12'h5A1;
20'b00000101100000100111 : ColourData = 12'h5A1;
20'b00000101110000100111 : ColourData = 12'h5A1;
20'b00000110000000100111 : ColourData = 12'h5A1;
20'b00000110010000100111 : ColourData = 12'h5A1;
20'b00000110100000100111 : ColourData = 12'h5A1;
20'b00000110110000100111 : ColourData = 12'h5A1;
20'b00000111000000100111 : ColourData = 12'h5A1;
20'b00000111010000100111 : ColourData = 12'h5A1;
20'b00000111100000100111 : ColourData = 12'h5A1;
20'b00000111110000100111 : ColourData = 12'h5A1;
20'b00001000000000100111 : ColourData = 12'h5A1;
20'b00001000010000100111 : ColourData = 12'h5A1;
20'b00001000100000100111 : ColourData = 12'h5A1;
20'b00001000110000100111 : ColourData = 12'h5A1;
20'b00001001000000100111 : ColourData = 12'h5A1;
20'b00001001010000100111 : ColourData = 12'h5A1;
20'b00001001100000100111 : ColourData = 12'h5A1;
20'b00001001110000100111 : ColourData = 12'h5A1;
20'b00001010000000100111 : ColourData = 12'h5A1;
20'b00001010010000100111 : ColourData = 12'h481;
20'b00001010100000100111 : ColourData = 12'h360;
20'b00001010110000100111 : ColourData = 12'h360;
20'b00001011000000100111 : ColourData = 12'h360;
20'b00001011010000100111 : ColourData = 12'h360;
20'b00001011100000100111 : ColourData = 12'h591;
20'b00001011110000100111 : ColourData = 12'h5A1;
20'b00001100000000100111 : ColourData = 12'h5A1;
20'b00001100010000100111 : ColourData = 12'h5A1;
20'b00001100100000100111 : ColourData = 12'h591;
20'b00001100110000100111 : ColourData = 12'h360;
20'b00001101000000100111 : ColourData = 12'h360;
20'b00001101010000100111 : ColourData = 12'h443;
20'b00001101100000100111 : ColourData = 12'h444;
20'b00001101110000100111 : ColourData = 12'h444;
20'b00001110000000100111 : ColourData = 12'h444;
20'b00001110010000100111 : ColourData = 12'h444;
20'b00001110100000100111 : ColourData = 12'h444;
20'b00001110110000100111 : ColourData = 12'h444;
20'b00000000000000101000 : ColourData = 12'h333;
20'b00000000010000101000 : ColourData = 12'h333;
20'b00000000100000101000 : ColourData = 12'h333;
20'b00000000110000101000 : ColourData = 12'h333;
20'b00000001000000101000 : ColourData = 12'h333;
20'b00000001010000101000 : ColourData = 12'h334;
20'b00000001100000101000 : ColourData = 12'h343;
20'b00000001110000101000 : ColourData = 12'h360;
20'b00000010000000101000 : ColourData = 12'h360;
20'b00000010010000101000 : ColourData = 12'h591;
20'b00000010100000101000 : ColourData = 12'h5A1;
20'b00000010110000101000 : ColourData = 12'h5A1;
20'b00000011000000101000 : ColourData = 12'h5A1;
20'b00000011010000101000 : ColourData = 12'h591;
20'b00000011100000101000 : ColourData = 12'h360;
20'b00000011110000101000 : ColourData = 12'h360;
20'b00000100000000101000 : ColourData = 12'h360;
20'b00000100010000101000 : ColourData = 12'h360;
20'b00000100100000101000 : ColourData = 12'h481;
20'b00000100110000101000 : ColourData = 12'h5A1;
20'b00000101000000101000 : ColourData = 12'h5A1;
20'b00000101010000101000 : ColourData = 12'h5A1;
20'b00000101100000101000 : ColourData = 12'h5A1;
20'b00000101110000101000 : ColourData = 12'h5A1;
20'b00000110000000101000 : ColourData = 12'h5A1;
20'b00000110010000101000 : ColourData = 12'h5A1;
20'b00000110100000101000 : ColourData = 12'h5A1;
20'b00000110110000101000 : ColourData = 12'h5A1;
20'b00000111000000101000 : ColourData = 12'h5A1;
20'b00000111010000101000 : ColourData = 12'h5A1;
20'b00000111100000101000 : ColourData = 12'h5A1;
20'b00000111110000101000 : ColourData = 12'h5A1;
20'b00001000000000101000 : ColourData = 12'h5A1;
20'b00001000010000101000 : ColourData = 12'h5A1;
20'b00001000100000101000 : ColourData = 12'h5A1;
20'b00001000110000101000 : ColourData = 12'h5A1;
20'b00001001000000101000 : ColourData = 12'h5A1;
20'b00001001010000101000 : ColourData = 12'h5A1;
20'b00001001100000101000 : ColourData = 12'h5A1;
20'b00001001110000101000 : ColourData = 12'h5A1;
20'b00001010000000101000 : ColourData = 12'h5A1;
20'b00001010010000101000 : ColourData = 12'h481;
20'b00001010100000101000 : ColourData = 12'h360;
20'b00001010110000101000 : ColourData = 12'h360;
20'b00001011000000101000 : ColourData = 12'h360;
20'b00001011010000101000 : ColourData = 12'h360;
20'b00001011100000101000 : ColourData = 12'h591;
20'b00001011110000101000 : ColourData = 12'h5A1;
20'b00001100000000101000 : ColourData = 12'h5A1;
20'b00001100010000101000 : ColourData = 12'h5A1;
20'b00001100100000101000 : ColourData = 12'h591;
20'b00001100110000101000 : ColourData = 12'h360;
20'b00001101000000101000 : ColourData = 12'h360;
20'b00001101010000101000 : ColourData = 12'h343;
20'b00001101100000101000 : ColourData = 12'h334;
20'b00001101110000101000 : ColourData = 12'h333;
20'b00001110000000101000 : ColourData = 12'h333;
20'b00001110010000101000 : ColourData = 12'h333;
20'b00001110100000101000 : ColourData = 12'h333;
20'b00001110110000101000 : ColourData = 12'h333;
20'b00000000000000101001 : ColourData = 12'h444;
20'b00000000010000101001 : ColourData = 12'h444;
20'b00000000100000101001 : ColourData = 12'h444;
20'b00000000110000101001 : ColourData = 12'h444;
20'b00000001000000101001 : ColourData = 12'h444;
20'b00000001010000101001 : ColourData = 12'h444;
20'b00000001100000101001 : ColourData = 12'h443;
20'b00000001110000101001 : ColourData = 12'h360;
20'b00000010000000101001 : ColourData = 12'h360;
20'b00000010010000101001 : ColourData = 12'h591;
20'b00000010100000101001 : ColourData = 12'h5A1;
20'b00000010110000101001 : ColourData = 12'h5A1;
20'b00000011000000101001 : ColourData = 12'h5A1;
20'b00000011010000101001 : ColourData = 12'h591;
20'b00000011100000101001 : ColourData = 12'h360;
20'b00000011110000101001 : ColourData = 12'h360;
20'b00000100000000101001 : ColourData = 12'h360;
20'b00000100010000101001 : ColourData = 12'h360;
20'b00000100100000101001 : ColourData = 12'h481;
20'b00000100110000101001 : ColourData = 12'h5A1;
20'b00000101000000101001 : ColourData = 12'h5A1;
20'b00000101010000101001 : ColourData = 12'h5A1;
20'b00000101100000101001 : ColourData = 12'h5A1;
20'b00000101110000101001 : ColourData = 12'h5A1;
20'b00000110000000101001 : ColourData = 12'h5A1;
20'b00000110010000101001 : ColourData = 12'h5A1;
20'b00000110100000101001 : ColourData = 12'h5A1;
20'b00000110110000101001 : ColourData = 12'h5A1;
20'b00000111000000101001 : ColourData = 12'h5A1;
20'b00000111010000101001 : ColourData = 12'h5A1;
20'b00000111100000101001 : ColourData = 12'h5A1;
20'b00000111110000101001 : ColourData = 12'h5A1;
20'b00001000000000101001 : ColourData = 12'h5A1;
20'b00001000010000101001 : ColourData = 12'h5A1;
20'b00001000100000101001 : ColourData = 12'h5A1;
20'b00001000110000101001 : ColourData = 12'h5A1;
20'b00001001000000101001 : ColourData = 12'h5A1;
20'b00001001010000101001 : ColourData = 12'h5A1;
20'b00001001100000101001 : ColourData = 12'h5A1;
20'b00001001110000101001 : ColourData = 12'h5A1;
20'b00001010000000101001 : ColourData = 12'h5A1;
20'b00001010010000101001 : ColourData = 12'h481;
20'b00001010100000101001 : ColourData = 12'h360;
20'b00001010110000101001 : ColourData = 12'h360;
20'b00001011000000101001 : ColourData = 12'h360;
20'b00001011010000101001 : ColourData = 12'h360;
20'b00001011100000101001 : ColourData = 12'h591;
20'b00001011110000101001 : ColourData = 12'h5A1;
20'b00001100000000101001 : ColourData = 12'h5A1;
20'b00001100010000101001 : ColourData = 12'h5A1;
20'b00001100100000101001 : ColourData = 12'h591;
20'b00001100110000101001 : ColourData = 12'h360;
20'b00001101000000101001 : ColourData = 12'h360;
20'b00001101010000101001 : ColourData = 12'h443;
20'b00001101100000101001 : ColourData = 12'h444;
20'b00001101110000101001 : ColourData = 12'h444;
20'b00001110000000101001 : ColourData = 12'h444;
20'b00001110010000101001 : ColourData = 12'h444;
20'b00001110100000101001 : ColourData = 12'h444;
20'b00001110110000101001 : ColourData = 12'h444;
20'b00000000000000101010 : ColourData = 12'h000;
20'b00000000010000101010 : ColourData = 12'h000;
20'b00000000100000101010 : ColourData = 12'h000;
20'b00000000110000101010 : ColourData = 12'h000;
20'b00000001000000101010 : ColourData = 12'h000;
20'b00000001010000101010 : ColourData = 12'h000;
20'b00000001100000101010 : ColourData = 12'h110;
20'b00000001110000101010 : ColourData = 12'h360;
20'b00000010000000101010 : ColourData = 12'h360;
20'b00000010010000101010 : ColourData = 12'h591;
20'b00000010100000101010 : ColourData = 12'h5A1;
20'b00000010110000101010 : ColourData = 12'h5A1;
20'b00000011000000101010 : ColourData = 12'h5A1;
20'b00000011010000101010 : ColourData = 12'h591;
20'b00000011100000101010 : ColourData = 12'h360;
20'b00000011110000101010 : ColourData = 12'h360;
20'b00000100000000101010 : ColourData = 12'h360;
20'b00000100010000101010 : ColourData = 12'h360;
20'b00000100100000101010 : ColourData = 12'h481;
20'b00000100110000101010 : ColourData = 12'h5A1;
20'b00000101000000101010 : ColourData = 12'h5A1;
20'b00000101010000101010 : ColourData = 12'h5A1;
20'b00000101100000101010 : ColourData = 12'h5A1;
20'b00000101110000101010 : ColourData = 12'h5A1;
20'b00000110000000101010 : ColourData = 12'h5A1;
20'b00000110010000101010 : ColourData = 12'h5A1;
20'b00000110100000101010 : ColourData = 12'h5A1;
20'b00000110110000101010 : ColourData = 12'h5A1;
20'b00000111000000101010 : ColourData = 12'h5A1;
20'b00000111010000101010 : ColourData = 12'h5A1;
20'b00000111100000101010 : ColourData = 12'h5A1;
20'b00000111110000101010 : ColourData = 12'h5A1;
20'b00001000000000101010 : ColourData = 12'h5A1;
20'b00001000010000101010 : ColourData = 12'h5A1;
20'b00001000100000101010 : ColourData = 12'h5A1;
20'b00001000110000101010 : ColourData = 12'h5A1;
20'b00001001000000101010 : ColourData = 12'h5A1;
20'b00001001010000101010 : ColourData = 12'h5A1;
20'b00001001100000101010 : ColourData = 12'h5A1;
20'b00001001110000101010 : ColourData = 12'h5A1;
20'b00001010000000101010 : ColourData = 12'h5A1;
20'b00001010010000101010 : ColourData = 12'h481;
20'b00001010100000101010 : ColourData = 12'h360;
20'b00001010110000101010 : ColourData = 12'h360;
20'b00001011000000101010 : ColourData = 12'h360;
20'b00001011010000101010 : ColourData = 12'h360;
20'b00001011100000101010 : ColourData = 12'h591;
20'b00001011110000101010 : ColourData = 12'h5A1;
20'b00001100000000101010 : ColourData = 12'h5A1;
20'b00001100010000101010 : ColourData = 12'h5A1;
20'b00001100100000101010 : ColourData = 12'h591;
20'b00001100110000101010 : ColourData = 12'h360;
20'b00001101000000101010 : ColourData = 12'h360;
20'b00001101010000101010 : ColourData = 12'h110;
20'b00001101100000101010 : ColourData = 12'h000;
20'b00001101110000101010 : ColourData = 12'h000;
20'b00001110000000101010 : ColourData = 12'h000;
20'b00001110010000101010 : ColourData = 12'h000;
20'b00001110100000101010 : ColourData = 12'h000;
20'b00001110110000101010 : ColourData = 12'h000;
20'b00000000000000101011 : ColourData = 12'h000;
20'b00000000010000101011 : ColourData = 12'h000;
20'b00000000100000101011 : ColourData = 12'h000;
20'b00000000110000101011 : ColourData = 12'h000;
20'b00000001000000101011 : ColourData = 12'h000;
20'b00000001010000101011 : ColourData = 12'h000;
20'b00000001100000101011 : ColourData = 12'h000;
20'b00000001110000101011 : ColourData = 12'h360;
20'b00000010000000101011 : ColourData = 12'h360;
20'b00000010010000101011 : ColourData = 12'h591;
20'b00000010100000101011 : ColourData = 12'h5A1;
20'b00000010110000101011 : ColourData = 12'h5A1;
20'b00000011000000101011 : ColourData = 12'h5A1;
20'b00000011010000101011 : ColourData = 12'h591;
20'b00000011100000101011 : ColourData = 12'h360;
20'b00000011110000101011 : ColourData = 12'h360;
20'b00000100000000101011 : ColourData = 12'h360;
20'b00000100010000101011 : ColourData = 12'h360;
20'b00000100100000101011 : ColourData = 12'h481;
20'b00000100110000101011 : ColourData = 12'h5A1;
20'b00000101000000101011 : ColourData = 12'h5A1;
20'b00000101010000101011 : ColourData = 12'h5A1;
20'b00000101100000101011 : ColourData = 12'h5A1;
20'b00000101110000101011 : ColourData = 12'h5A1;
20'b00000110000000101011 : ColourData = 12'h5A1;
20'b00000110010000101011 : ColourData = 12'h5A1;
20'b00000110100000101011 : ColourData = 12'h5A1;
20'b00000110110000101011 : ColourData = 12'h5A1;
20'b00000111000000101011 : ColourData = 12'h5A1;
20'b00000111010000101011 : ColourData = 12'h5A1;
20'b00000111100000101011 : ColourData = 12'h5A1;
20'b00000111110000101011 : ColourData = 12'h5A1;
20'b00001000000000101011 : ColourData = 12'h5A1;
20'b00001000010000101011 : ColourData = 12'h5A1;
20'b00001000100000101011 : ColourData = 12'h5A1;
20'b00001000110000101011 : ColourData = 12'h5A1;
20'b00001001000000101011 : ColourData = 12'h5A1;
20'b00001001010000101011 : ColourData = 12'h5A1;
20'b00001001100000101011 : ColourData = 12'h5A1;
20'b00001001110000101011 : ColourData = 12'h5A1;
20'b00001010000000101011 : ColourData = 12'h5A1;
20'b00001010010000101011 : ColourData = 12'h481;
20'b00001010100000101011 : ColourData = 12'h360;
20'b00001010110000101011 : ColourData = 12'h360;
20'b00001011000000101011 : ColourData = 12'h360;
20'b00001011010000101011 : ColourData = 12'h360;
20'b00001011100000101011 : ColourData = 12'h591;
20'b00001011110000101011 : ColourData = 12'h5A1;
20'b00001100000000101011 : ColourData = 12'h5A1;
20'b00001100010000101011 : ColourData = 12'h5A1;
20'b00001100100000101011 : ColourData = 12'h591;
20'b00001100110000101011 : ColourData = 12'h360;
20'b00001101000000101011 : ColourData = 12'h360;
20'b00001101010000101011 : ColourData = 12'h000;
20'b00001101100000101011 : ColourData = 12'h000;
20'b00001101110000101011 : ColourData = 12'h000;
20'b00001110000000101011 : ColourData = 12'h000;
20'b00001110010000101011 : ColourData = 12'h000;
20'b00001110100000101011 : ColourData = 12'h000;
20'b00001110110000101011 : ColourData = 12'h000;
20'b00000000000000101100 : ColourData = 12'h333;
20'b00000000010000101100 : ColourData = 12'h333;
20'b00000000100000101100 : ColourData = 12'h333;
20'b00000000110000101100 : ColourData = 12'h333;
20'b00000001000000101100 : ColourData = 12'h333;
20'b00000001010000101100 : ColourData = 12'h333;
20'b00000001100000101100 : ColourData = 12'h333;
20'b00000001110000101100 : ColourData = 12'h360;
20'b00000010000000101100 : ColourData = 12'h360;
20'b00000010010000101100 : ColourData = 12'h591;
20'b00000010100000101100 : ColourData = 12'h5A1;
20'b00000010110000101100 : ColourData = 12'h5A1;
20'b00000011000000101100 : ColourData = 12'h5A1;
20'b00000011010000101100 : ColourData = 12'h591;
20'b00000011100000101100 : ColourData = 12'h360;
20'b00000011110000101100 : ColourData = 12'h360;
20'b00000100000000101100 : ColourData = 12'h360;
20'b00000100010000101100 : ColourData = 12'h360;
20'b00000100100000101100 : ColourData = 12'h481;
20'b00000100110000101100 : ColourData = 12'h5A1;
20'b00000101000000101100 : ColourData = 12'h5A1;
20'b00000101010000101100 : ColourData = 12'h5A1;
20'b00000101100000101100 : ColourData = 12'h5A1;
20'b00000101110000101100 : ColourData = 12'h5A1;
20'b00000110000000101100 : ColourData = 12'h5A1;
20'b00000110010000101100 : ColourData = 12'h5A1;
20'b00000110100000101100 : ColourData = 12'h5A1;
20'b00000110110000101100 : ColourData = 12'h5A1;
20'b00000111000000101100 : ColourData = 12'h5A1;
20'b00000111010000101100 : ColourData = 12'h5A1;
20'b00000111100000101100 : ColourData = 12'h5A1;
20'b00000111110000101100 : ColourData = 12'h5A1;
20'b00001000000000101100 : ColourData = 12'h5A1;
20'b00001000010000101100 : ColourData = 12'h5A1;
20'b00001000100000101100 : ColourData = 12'h5A1;
20'b00001000110000101100 : ColourData = 12'h5A1;
20'b00001001000000101100 : ColourData = 12'h5A1;
20'b00001001010000101100 : ColourData = 12'h5A1;
20'b00001001100000101100 : ColourData = 12'h5A1;
20'b00001001110000101100 : ColourData = 12'h5A1;
20'b00001010000000101100 : ColourData = 12'h5A1;
20'b00001010010000101100 : ColourData = 12'h481;
20'b00001010100000101100 : ColourData = 12'h360;
20'b00001010110000101100 : ColourData = 12'h360;
20'b00001011000000101100 : ColourData = 12'h360;
20'b00001011010000101100 : ColourData = 12'h360;
20'b00001011100000101100 : ColourData = 12'h591;
20'b00001011110000101100 : ColourData = 12'h5A1;
20'b00001100000000101100 : ColourData = 12'h5A1;
20'b00001100010000101100 : ColourData = 12'h5A1;
20'b00001100100000101100 : ColourData = 12'h591;
20'b00001100110000101100 : ColourData = 12'h360;
20'b00001101000000101100 : ColourData = 12'h360;
20'b00001101010000101100 : ColourData = 12'h333;
20'b00001101100000101100 : ColourData = 12'h333;
20'b00001101110000101100 : ColourData = 12'h333;
20'b00001110000000101100 : ColourData = 12'h333;
20'b00001110010000101100 : ColourData = 12'h333;
20'b00001110100000101100 : ColourData = 12'h333;
20'b00001110110000101100 : ColourData = 12'h333;
20'b00000000000000101101 : ColourData = 12'h333;
20'b00000000010000101101 : ColourData = 12'h333;
20'b00000000100000101101 : ColourData = 12'h333;
20'b00000000110000101101 : ColourData = 12'h333;
20'b00000001000000101101 : ColourData = 12'h333;
20'b00000001010000101101 : ColourData = 12'h333;
20'b00000001100000101101 : ColourData = 12'h333;
20'b00000001110000101101 : ColourData = 12'h360;
20'b00000010000000101101 : ColourData = 12'h360;
20'b00000010010000101101 : ColourData = 12'h591;
20'b00000010100000101101 : ColourData = 12'h5A1;
20'b00000010110000101101 : ColourData = 12'h5A1;
20'b00000011000000101101 : ColourData = 12'h5A1;
20'b00000011010000101101 : ColourData = 12'h591;
20'b00000011100000101101 : ColourData = 12'h360;
20'b00000011110000101101 : ColourData = 12'h360;
20'b00000100000000101101 : ColourData = 12'h360;
20'b00000100010000101101 : ColourData = 12'h360;
20'b00000100100000101101 : ColourData = 12'h481;
20'b00000100110000101101 : ColourData = 12'h5A1;
20'b00000101000000101101 : ColourData = 12'h5A1;
20'b00000101010000101101 : ColourData = 12'h5A1;
20'b00000101100000101101 : ColourData = 12'h5A1;
20'b00000101110000101101 : ColourData = 12'h5A1;
20'b00000110000000101101 : ColourData = 12'h5A1;
20'b00000110010000101101 : ColourData = 12'h5A1;
20'b00000110100000101101 : ColourData = 12'h5A1;
20'b00000110110000101101 : ColourData = 12'h5A1;
20'b00000111000000101101 : ColourData = 12'h5A1;
20'b00000111010000101101 : ColourData = 12'h5A1;
20'b00000111100000101101 : ColourData = 12'h5A1;
20'b00000111110000101101 : ColourData = 12'h5A1;
20'b00001000000000101101 : ColourData = 12'h5A1;
20'b00001000010000101101 : ColourData = 12'h5A1;
20'b00001000100000101101 : ColourData = 12'h5A1;
20'b00001000110000101101 : ColourData = 12'h5A1;
20'b00001001000000101101 : ColourData = 12'h5A1;
20'b00001001010000101101 : ColourData = 12'h5A1;
20'b00001001100000101101 : ColourData = 12'h5A1;
20'b00001001110000101101 : ColourData = 12'h5A1;
20'b00001010000000101101 : ColourData = 12'h5A1;
20'b00001010010000101101 : ColourData = 12'h481;
20'b00001010100000101101 : ColourData = 12'h360;
20'b00001010110000101101 : ColourData = 12'h360;
20'b00001011000000101101 : ColourData = 12'h360;
20'b00001011010000101101 : ColourData = 12'h360;
20'b00001011100000101101 : ColourData = 12'h591;
20'b00001011110000101101 : ColourData = 12'h5A1;
20'b00001100000000101101 : ColourData = 12'h5A1;
20'b00001100010000101101 : ColourData = 12'h5A1;
20'b00001100100000101101 : ColourData = 12'h591;
20'b00001100110000101101 : ColourData = 12'h360;
20'b00001101000000101101 : ColourData = 12'h360;
20'b00001101010000101101 : ColourData = 12'h333;
20'b00001101100000101101 : ColourData = 12'h333;
20'b00001101110000101101 : ColourData = 12'h333;
20'b00001110000000101101 : ColourData = 12'h333;
20'b00001110010000101101 : ColourData = 12'h333;
20'b00001110100000101101 : ColourData = 12'h333;
20'b00001110110000101101 : ColourData = 12'h333;
20'b00000000000000101110 : ColourData = 12'h000;
20'b00000000010000101110 : ColourData = 12'h000;
20'b00000000100000101110 : ColourData = 12'h000;
20'b00000000110000101110 : ColourData = 12'h000;
20'b00000001000000101110 : ColourData = 12'h000;
20'b00000001010000101110 : ColourData = 12'h000;
20'b00000001100000101110 : ColourData = 12'h000;
20'b00000001110000101110 : ColourData = 12'h360;
20'b00000010000000101110 : ColourData = 12'h360;
20'b00000010010000101110 : ColourData = 12'h591;
20'b00000010100000101110 : ColourData = 12'h5A1;
20'b00000010110000101110 : ColourData = 12'h5A1;
20'b00000011000000101110 : ColourData = 12'h5A1;
20'b00000011010000101110 : ColourData = 12'h591;
20'b00000011100000101110 : ColourData = 12'h360;
20'b00000011110000101110 : ColourData = 12'h360;
20'b00000100000000101110 : ColourData = 12'h360;
20'b00000100010000101110 : ColourData = 12'h360;
20'b00000100100000101110 : ColourData = 12'h481;
20'b00000100110000101110 : ColourData = 12'h6A1;
20'b00000101000000101110 : ColourData = 12'h5A1;
20'b00000101010000101110 : ColourData = 12'h5A1;
20'b00000101100000101110 : ColourData = 12'h5A1;
20'b00000101110000101110 : ColourData = 12'h5A1;
20'b00000110000000101110 : ColourData = 12'h5A1;
20'b00000110010000101110 : ColourData = 12'h5A1;
20'b00000110100000101110 : ColourData = 12'h5A1;
20'b00000110110000101110 : ColourData = 12'h5A1;
20'b00000111000000101110 : ColourData = 12'h5A1;
20'b00000111010000101110 : ColourData = 12'h5A1;
20'b00000111100000101110 : ColourData = 12'h5A1;
20'b00000111110000101110 : ColourData = 12'h5A1;
20'b00001000000000101110 : ColourData = 12'h5A1;
20'b00001000010000101110 : ColourData = 12'h5A1;
20'b00001000100000101110 : ColourData = 12'h5A1;
20'b00001000110000101110 : ColourData = 12'h5A1;
20'b00001001000000101110 : ColourData = 12'h5A1;
20'b00001001010000101110 : ColourData = 12'h5A1;
20'b00001001100000101110 : ColourData = 12'h5A1;
20'b00001001110000101110 : ColourData = 12'h5A1;
20'b00001010000000101110 : ColourData = 12'h6A1;
20'b00001010010000101110 : ColourData = 12'h481;
20'b00001010100000101110 : ColourData = 12'h360;
20'b00001010110000101110 : ColourData = 12'h360;
20'b00001011000000101110 : ColourData = 12'h360;
20'b00001011010000101110 : ColourData = 12'h360;
20'b00001011100000101110 : ColourData = 12'h591;
20'b00001011110000101110 : ColourData = 12'h5A1;
20'b00001100000000101110 : ColourData = 12'h5A1;
20'b00001100010000101110 : ColourData = 12'h5A1;
20'b00001100100000101110 : ColourData = 12'h591;
20'b00001100110000101110 : ColourData = 12'h360;
20'b00001101000000101110 : ColourData = 12'h360;
20'b00001101010000101110 : ColourData = 12'h000;
20'b00001101100000101110 : ColourData = 12'h000;
20'b00001101110000101110 : ColourData = 12'h000;
20'b00001110000000101110 : ColourData = 12'h000;
20'b00001110010000101110 : ColourData = 12'h000;
20'b00001110100000101110 : ColourData = 12'h000;
20'b00001110110000101110 : ColourData = 12'h000;
20'b00000000000000101111 : ColourData = 12'h000;
20'b00000000010000101111 : ColourData = 12'h000;
20'b00000000100000101111 : ColourData = 12'h000;
20'b00000000110000101111 : ColourData = 12'h000;
20'b00000001000000101111 : ColourData = 12'h000;
20'b00000001010000101111 : ColourData = 12'h000;
20'b00000001100000101111 : ColourData = 12'h110;
20'b00000001110000101111 : ColourData = 12'h360;
20'b00000010000000101111 : ColourData = 12'h360;
20'b00000010010000101111 : ColourData = 12'h591;
20'b00000010100000101111 : ColourData = 12'h5A1;
20'b00000010110000101111 : ColourData = 12'h5A1;
20'b00000011000000101111 : ColourData = 12'h5A1;
20'b00000011010000101111 : ColourData = 12'h591;
20'b00000011100000101111 : ColourData = 12'h360;
20'b00000011110000101111 : ColourData = 12'h360;
20'b00000100000000101111 : ColourData = 12'h360;
20'b00000100010000101111 : ColourData = 12'h360;
20'b00000100100000101111 : ColourData = 12'h471;
20'b00000100110000101111 : ColourData = 12'h591;
20'b00000101000000101111 : ColourData = 12'h581;
20'b00000101010000101111 : ColourData = 12'h581;
20'b00000101100000101111 : ColourData = 12'h581;
20'b00000101110000101111 : ColourData = 12'h581;
20'b00000110000000101111 : ColourData = 12'h581;
20'b00000110010000101111 : ColourData = 12'h581;
20'b00000110100000101111 : ColourData = 12'h581;
20'b00000110110000101111 : ColourData = 12'h581;
20'b00000111000000101111 : ColourData = 12'h581;
20'b00000111010000101111 : ColourData = 12'h581;
20'b00000111100000101111 : ColourData = 12'h581;
20'b00000111110000101111 : ColourData = 12'h581;
20'b00001000000000101111 : ColourData = 12'h581;
20'b00001000010000101111 : ColourData = 12'h581;
20'b00001000100000101111 : ColourData = 12'h581;
20'b00001000110000101111 : ColourData = 12'h581;
20'b00001001000000101111 : ColourData = 12'h581;
20'b00001001010000101111 : ColourData = 12'h581;
20'b00001001100000101111 : ColourData = 12'h581;
20'b00001001110000101111 : ColourData = 12'h581;
20'b00001010000000101111 : ColourData = 12'h591;
20'b00001010010000101111 : ColourData = 12'h471;
20'b00001010100000101111 : ColourData = 12'h360;
20'b00001010110000101111 : ColourData = 12'h360;
20'b00001011000000101111 : ColourData = 12'h360;
20'b00001011010000101111 : ColourData = 12'h360;
20'b00001011100000101111 : ColourData = 12'h591;
20'b00001011110000101111 : ColourData = 12'h5A1;
20'b00001100000000101111 : ColourData = 12'h5A1;
20'b00001100010000101111 : ColourData = 12'h5A1;
20'b00001100100000101111 : ColourData = 12'h591;
20'b00001100110000101111 : ColourData = 12'h360;
20'b00001101000000101111 : ColourData = 12'h360;
20'b00001101010000101111 : ColourData = 12'h110;
20'b00001101100000101111 : ColourData = 12'h000;
20'b00001101110000101111 : ColourData = 12'h000;
20'b00001110000000101111 : ColourData = 12'h000;
20'b00001110010000101111 : ColourData = 12'h000;
20'b00001110100000101111 : ColourData = 12'h000;
20'b00001110110000101111 : ColourData = 12'h000;
20'b00000000000000110000 : ColourData = 12'h444;
20'b00000000010000110000 : ColourData = 12'h444;
20'b00000000100000110000 : ColourData = 12'h444;
20'b00000000110000110000 : ColourData = 12'h444;
20'b00000001000000110000 : ColourData = 12'h444;
20'b00000001010000110000 : ColourData = 12'h444;
20'b00000001100000110000 : ColourData = 12'h444;
20'b00000001110000110000 : ColourData = 12'h360;
20'b00000010000000110000 : ColourData = 12'h360;
20'b00000010010000110000 : ColourData = 12'h591;
20'b00000010100000110000 : ColourData = 12'h5A1;
20'b00000010110000110000 : ColourData = 12'h5A1;
20'b00000011000000110000 : ColourData = 12'h5A1;
20'b00000011010000110000 : ColourData = 12'h591;
20'b00000011100000110000 : ColourData = 12'h360;
20'b00000011110000110000 : ColourData = 12'h360;
20'b00000100000000110000 : ColourData = 12'h360;
20'b00000100010000110000 : ColourData = 12'h360;
20'b00000100100000110000 : ColourData = 12'h360;
20'b00000100110000110000 : ColourData = 12'h360;
20'b00000101000000110000 : ColourData = 12'h360;
20'b00000101010000110000 : ColourData = 12'h360;
20'b00000101100000110000 : ColourData = 12'h360;
20'b00000101110000110000 : ColourData = 12'h360;
20'b00000110000000110000 : ColourData = 12'h360;
20'b00000110010000110000 : ColourData = 12'h360;
20'b00000110100000110000 : ColourData = 12'h360;
20'b00000110110000110000 : ColourData = 12'h360;
20'b00000111000000110000 : ColourData = 12'h360;
20'b00000111010000110000 : ColourData = 12'h360;
20'b00000111100000110000 : ColourData = 12'h360;
20'b00000111110000110000 : ColourData = 12'h360;
20'b00001000000000110000 : ColourData = 12'h360;
20'b00001000010000110000 : ColourData = 12'h360;
20'b00001000100000110000 : ColourData = 12'h360;
20'b00001000110000110000 : ColourData = 12'h360;
20'b00001001000000110000 : ColourData = 12'h360;
20'b00001001010000110000 : ColourData = 12'h360;
20'b00001001100000110000 : ColourData = 12'h360;
20'b00001001110000110000 : ColourData = 12'h360;
20'b00001010000000110000 : ColourData = 12'h360;
20'b00001010010000110000 : ColourData = 12'h360;
20'b00001010100000110000 : ColourData = 12'h360;
20'b00001010110000110000 : ColourData = 12'h360;
20'b00001011000000110000 : ColourData = 12'h360;
20'b00001011010000110000 : ColourData = 12'h360;
20'b00001011100000110000 : ColourData = 12'h591;
20'b00001011110000110000 : ColourData = 12'h5A1;
20'b00001100000000110000 : ColourData = 12'h5A1;
20'b00001100010000110000 : ColourData = 12'h5A1;
20'b00001100100000110000 : ColourData = 12'h591;
20'b00001100110000110000 : ColourData = 12'h360;
20'b00001101000000110000 : ColourData = 12'h360;
20'b00001101010000110000 : ColourData = 12'h444;
20'b00001101100000110000 : ColourData = 12'h444;
20'b00001101110000110000 : ColourData = 12'h444;
20'b00001110000000110000 : ColourData = 12'h444;
20'b00001110010000110000 : ColourData = 12'h444;
20'b00001110100000110000 : ColourData = 12'h444;
20'b00001110110000110000 : ColourData = 12'h444;
20'b00000000000000110001 : ColourData = 12'h111;
20'b00000000010000110001 : ColourData = 12'h111;
20'b00000000100000110001 : ColourData = 12'h111;
20'b00000000110000110001 : ColourData = 12'h111;
20'b00000001000000110001 : ColourData = 12'h111;
20'b00000001010000110001 : ColourData = 12'h111;
20'b00000001100000110001 : ColourData = 12'h111;
20'b00000001110000110001 : ColourData = 12'h360;
20'b00000010000000110001 : ColourData = 12'h360;
20'b00000010010000110001 : ColourData = 12'h591;
20'b00000010100000110001 : ColourData = 12'h5A1;
20'b00000010110000110001 : ColourData = 12'h5A1;
20'b00000011000000110001 : ColourData = 12'h5A1;
20'b00000011010000110001 : ColourData = 12'h591;
20'b00000011100000110001 : ColourData = 12'h481;
20'b00000011110000110001 : ColourData = 12'h481;
20'b00000100000000110001 : ColourData = 12'h360;
20'b00000100010000110001 : ColourData = 12'h360;
20'b00000100100000110001 : ColourData = 12'h360;
20'b00000100110000110001 : ColourData = 12'h360;
20'b00000101000000110001 : ColourData = 12'h360;
20'b00000101010000110001 : ColourData = 12'h360;
20'b00000101100000110001 : ColourData = 12'h360;
20'b00000101110000110001 : ColourData = 12'h360;
20'b00000110000000110001 : ColourData = 12'h360;
20'b00000110010000110001 : ColourData = 12'h360;
20'b00000110100000110001 : ColourData = 12'h360;
20'b00000110110000110001 : ColourData = 12'h360;
20'b00000111000000110001 : ColourData = 12'h360;
20'b00000111010000110001 : ColourData = 12'h360;
20'b00000111100000110001 : ColourData = 12'h360;
20'b00000111110000110001 : ColourData = 12'h360;
20'b00001000000000110001 : ColourData = 12'h360;
20'b00001000010000110001 : ColourData = 12'h360;
20'b00001000100000110001 : ColourData = 12'h360;
20'b00001000110000110001 : ColourData = 12'h360;
20'b00001001000000110001 : ColourData = 12'h360;
20'b00001001010000110001 : ColourData = 12'h360;
20'b00001001100000110001 : ColourData = 12'h360;
20'b00001001110000110001 : ColourData = 12'h360;
20'b00001010000000110001 : ColourData = 12'h360;
20'b00001010010000110001 : ColourData = 12'h360;
20'b00001010100000110001 : ColourData = 12'h360;
20'b00001010110000110001 : ColourData = 12'h360;
20'b00001011000000110001 : ColourData = 12'h481;
20'b00001011010000110001 : ColourData = 12'h481;
20'b00001011100000110001 : ColourData = 12'h591;
20'b00001011110000110001 : ColourData = 12'h5A1;
20'b00001100000000110001 : ColourData = 12'h5A1;
20'b00001100010000110001 : ColourData = 12'h5A1;
20'b00001100100000110001 : ColourData = 12'h591;
20'b00001100110000110001 : ColourData = 12'h360;
20'b00001101000000110001 : ColourData = 12'h360;
20'b00001101010000110001 : ColourData = 12'h111;
20'b00001101100000110001 : ColourData = 12'h111;
20'b00001101110000110001 : ColourData = 12'h111;
20'b00001110000000110001 : ColourData = 12'h111;
20'b00001110010000110001 : ColourData = 12'h111;
20'b00001110100000110001 : ColourData = 12'h111;
20'b00001110110000110001 : ColourData = 12'h111;
20'b00000000000000110010 : ColourData = 12'h000;
20'b00000000010000110010 : ColourData = 12'h000;
20'b00000000100000110010 : ColourData = 12'h000;
20'b00000000110000110010 : ColourData = 12'h000;
20'b00000001000000110010 : ColourData = 12'h000;
20'b00000001010000110010 : ColourData = 12'h000;
20'b00000001100000110010 : ColourData = 12'h000;
20'b00000001110000110010 : ColourData = 12'h360;
20'b00000010000000110010 : ColourData = 12'h360;
20'b00000010010000110010 : ColourData = 12'h591;
20'b00000010100000110010 : ColourData = 12'h5A1;
20'b00000010110000110010 : ColourData = 12'h5A1;
20'b00000011000000110010 : ColourData = 12'h5A1;
20'b00000011010000110010 : ColourData = 12'h5A1;
20'b00000011100000110010 : ColourData = 12'h5A1;
20'b00000011110000110010 : ColourData = 12'h5A1;
20'b00000100000000110010 : ColourData = 12'h360;
20'b00000100010000110010 : ColourData = 12'h360;
20'b00000100100000110010 : ColourData = 12'h360;
20'b00000100110000110010 : ColourData = 12'h360;
20'b00000101000000110010 : ColourData = 12'h360;
20'b00000101010000110010 : ColourData = 12'h360;
20'b00000101100000110010 : ColourData = 12'h360;
20'b00000101110000110010 : ColourData = 12'h360;
20'b00000110000000110010 : ColourData = 12'h360;
20'b00000110010000110010 : ColourData = 12'h360;
20'b00000110100000110010 : ColourData = 12'h360;
20'b00000110110000110010 : ColourData = 12'h360;
20'b00000111000000110010 : ColourData = 12'h360;
20'b00000111010000110010 : ColourData = 12'h360;
20'b00000111100000110010 : ColourData = 12'h360;
20'b00000111110000110010 : ColourData = 12'h360;
20'b00001000000000110010 : ColourData = 12'h360;
20'b00001000010000110010 : ColourData = 12'h360;
20'b00001000100000110010 : ColourData = 12'h360;
20'b00001000110000110010 : ColourData = 12'h360;
20'b00001001000000110010 : ColourData = 12'h360;
20'b00001001010000110010 : ColourData = 12'h360;
20'b00001001100000110010 : ColourData = 12'h360;
20'b00001001110000110010 : ColourData = 12'h360;
20'b00001010000000110010 : ColourData = 12'h360;
20'b00001010010000110010 : ColourData = 12'h360;
20'b00001010100000110010 : ColourData = 12'h360;
20'b00001010110000110010 : ColourData = 12'h360;
20'b00001011000000110010 : ColourData = 12'h5A1;
20'b00001011010000110010 : ColourData = 12'h5A1;
20'b00001011100000110010 : ColourData = 12'h5A1;
20'b00001011110000110010 : ColourData = 12'h5A1;
20'b00001100000000110010 : ColourData = 12'h5A1;
20'b00001100010000110010 : ColourData = 12'h5A1;
20'b00001100100000110010 : ColourData = 12'h591;
20'b00001100110000110010 : ColourData = 12'h360;
20'b00001101000000110010 : ColourData = 12'h360;
20'b00001101010000110010 : ColourData = 12'h000;
20'b00001101100000110010 : ColourData = 12'h000;
20'b00001101110000110010 : ColourData = 12'h000;
20'b00001110000000110010 : ColourData = 12'h000;
20'b00001110010000110010 : ColourData = 12'h000;
20'b00001110100000110010 : ColourData = 12'h000;
20'b00001110110000110010 : ColourData = 12'h000;
20'b00000000000000110011 : ColourData = 12'h333;
20'b00000000010000110011 : ColourData = 12'h333;
20'b00000000100000110011 : ColourData = 12'h333;
20'b00000000110000110011 : ColourData = 12'h333;
20'b00000001000000110011 : ColourData = 12'h333;
20'b00000001010000110011 : ColourData = 12'h333;
20'b00000001100000110011 : ColourData = 12'h333;
20'b00000001110000110011 : ColourData = 12'h360;
20'b00000010000000110011 : ColourData = 12'h360;
20'b00000010010000110011 : ColourData = 12'h591;
20'b00000010100000110011 : ColourData = 12'h5A1;
20'b00000010110000110011 : ColourData = 12'h5A1;
20'b00000011000000110011 : ColourData = 12'h5A1;
20'b00000011010000110011 : ColourData = 12'h5A1;
20'b00000011100000110011 : ColourData = 12'h5A1;
20'b00000011110000110011 : ColourData = 12'h5A1;
20'b00000100000000110011 : ColourData = 12'h591;
20'b00000100010000110011 : ColourData = 12'h591;
20'b00000100100000110011 : ColourData = 12'h591;
20'b00000100110000110011 : ColourData = 12'h591;
20'b00000101000000110011 : ColourData = 12'h591;
20'b00000101010000110011 : ColourData = 12'h591;
20'b00000101100000110011 : ColourData = 12'h591;
20'b00000101110000110011 : ColourData = 12'h591;
20'b00000110000000110011 : ColourData = 12'h591;
20'b00000110010000110011 : ColourData = 12'h591;
20'b00000110100000110011 : ColourData = 12'h591;
20'b00000110110000110011 : ColourData = 12'h481;
20'b00000111000000110011 : ColourData = 12'h360;
20'b00000111010000110011 : ColourData = 12'h360;
20'b00000111100000110011 : ColourData = 12'h360;
20'b00000111110000110011 : ColourData = 12'h360;
20'b00001000000000110011 : ColourData = 12'h481;
20'b00001000010000110011 : ColourData = 12'h591;
20'b00001000100000110011 : ColourData = 12'h591;
20'b00001000110000110011 : ColourData = 12'h591;
20'b00001001000000110011 : ColourData = 12'h591;
20'b00001001010000110011 : ColourData = 12'h591;
20'b00001001100000110011 : ColourData = 12'h591;
20'b00001001110000110011 : ColourData = 12'h591;
20'b00001010000000110011 : ColourData = 12'h591;
20'b00001010010000110011 : ColourData = 12'h591;
20'b00001010100000110011 : ColourData = 12'h591;
20'b00001010110000110011 : ColourData = 12'h591;
20'b00001011000000110011 : ColourData = 12'h5A1;
20'b00001011010000110011 : ColourData = 12'h5A1;
20'b00001011100000110011 : ColourData = 12'h5A1;
20'b00001011110000110011 : ColourData = 12'h5A1;
20'b00001100000000110011 : ColourData = 12'h5A1;
20'b00001100010000110011 : ColourData = 12'h5A1;
20'b00001100100000110011 : ColourData = 12'h591;
20'b00001100110000110011 : ColourData = 12'h360;
20'b00001101000000110011 : ColourData = 12'h360;
20'b00001101010000110011 : ColourData = 12'h333;
20'b00001101100000110011 : ColourData = 12'h333;
20'b00001101110000110011 : ColourData = 12'h333;
20'b00001110000000110011 : ColourData = 12'h333;
20'b00001110010000110011 : ColourData = 12'h333;
20'b00001110100000110011 : ColourData = 12'h333;
20'b00001110110000110011 : ColourData = 12'h333;
20'b00000000000000110100 : ColourData = 12'h333;
20'b00000000010000110100 : ColourData = 12'h333;
20'b00000000100000110100 : ColourData = 12'h333;
20'b00000000110000110100 : ColourData = 12'h333;
20'b00000001000000110100 : ColourData = 12'h333;
20'b00000001010000110100 : ColourData = 12'h333;
20'b00000001100000110100 : ColourData = 12'h343;
20'b00000001110000110100 : ColourData = 12'h360;
20'b00000010000000110100 : ColourData = 12'h360;
20'b00000010010000110100 : ColourData = 12'h591;
20'b00000010100000110100 : ColourData = 12'h591;
20'b00000010110000110100 : ColourData = 12'h591;
20'b00000011000000110100 : ColourData = 12'h5A1;
20'b00000011010000110100 : ColourData = 12'h5A1;
20'b00000011100000110100 : ColourData = 12'h5A1;
20'b00000011110000110100 : ColourData = 12'h5A1;
20'b00000100000000110100 : ColourData = 12'h5A1;
20'b00000100010000110100 : ColourData = 12'h5A1;
20'b00000100100000110100 : ColourData = 12'h5A1;
20'b00000100110000110100 : ColourData = 12'h5A1;
20'b00000101000000110100 : ColourData = 12'h5A1;
20'b00000101010000110100 : ColourData = 12'h5A1;
20'b00000101100000110100 : ColourData = 12'h5A1;
20'b00000101110000110100 : ColourData = 12'h5A1;
20'b00000110000000110100 : ColourData = 12'h5A1;
20'b00000110010000110100 : ColourData = 12'h5A1;
20'b00000110100000110100 : ColourData = 12'h5A1;
20'b00000110110000110100 : ColourData = 12'h591;
20'b00000111000000110100 : ColourData = 12'h360;
20'b00000111010000110100 : ColourData = 12'h360;
20'b00000111100000110100 : ColourData = 12'h360;
20'b00000111110000110100 : ColourData = 12'h360;
20'b00001000000000110100 : ColourData = 12'h591;
20'b00001000010000110100 : ColourData = 12'h5A1;
20'b00001000100000110100 : ColourData = 12'h5A1;
20'b00001000110000110100 : ColourData = 12'h5A1;
20'b00001001000000110100 : ColourData = 12'h5A1;
20'b00001001010000110100 : ColourData = 12'h5A1;
20'b00001001100000110100 : ColourData = 12'h5A1;
20'b00001001110000110100 : ColourData = 12'h5A1;
20'b00001010000000110100 : ColourData = 12'h5A1;
20'b00001010010000110100 : ColourData = 12'h5A1;
20'b00001010100000110100 : ColourData = 12'h5A1;
20'b00001010110000110100 : ColourData = 12'h5A1;
20'b00001011000000110100 : ColourData = 12'h5A1;
20'b00001011010000110100 : ColourData = 12'h5A1;
20'b00001011100000110100 : ColourData = 12'h5A1;
20'b00001011110000110100 : ColourData = 12'h5A1;
20'b00001100000000110100 : ColourData = 12'h591;
20'b00001100010000110100 : ColourData = 12'h591;
20'b00001100100000110100 : ColourData = 12'h591;
20'b00001100110000110100 : ColourData = 12'h360;
20'b00001101000000110100 : ColourData = 12'h360;
20'b00001101010000110100 : ColourData = 12'h343;
20'b00001101100000110100 : ColourData = 12'h333;
20'b00001101110000110100 : ColourData = 12'h333;
20'b00001110000000110100 : ColourData = 12'h333;
20'b00001110010000110100 : ColourData = 12'h333;
20'b00001110100000110100 : ColourData = 12'h333;
20'b00001110110000110100 : ColourData = 12'h333;
20'b00000000000000110101 : ColourData = 12'h000;
20'b00000000010000110101 : ColourData = 12'h000;
20'b00000000100000110101 : ColourData = 12'h000;
20'b00000000110000110101 : ColourData = 12'h000;
20'b00000001000000110101 : ColourData = 12'h000;
20'b00000001010000110101 : ColourData = 12'h000;
20'b00000001100000110101 : ColourData = 12'h000;
20'b00000001110000110101 : ColourData = 12'h360;
20'b00000010000000110101 : ColourData = 12'h360;
20'b00000010010000110101 : ColourData = 12'h360;
20'b00000010100000110101 : ColourData = 12'h360;
20'b00000010110000110101 : ColourData = 12'h481;
20'b00000011000000110101 : ColourData = 12'h6A1;
20'b00000011010000110101 : ColourData = 12'h5A1;
20'b00000011100000110101 : ColourData = 12'h5A1;
20'b00000011110000110101 : ColourData = 12'h5A1;
20'b00000100000000110101 : ColourData = 12'h5A1;
20'b00000100010000110101 : ColourData = 12'h5A1;
20'b00000100100000110101 : ColourData = 12'h5A1;
20'b00000100110000110101 : ColourData = 12'h5A1;
20'b00000101000000110101 : ColourData = 12'h5A1;
20'b00000101010000110101 : ColourData = 12'h5A1;
20'b00000101100000110101 : ColourData = 12'h5A1;
20'b00000101110000110101 : ColourData = 12'h5A1;
20'b00000110000000110101 : ColourData = 12'h5A1;
20'b00000110010000110101 : ColourData = 12'h5A1;
20'b00000110100000110101 : ColourData = 12'h5A1;
20'b00000110110000110101 : ColourData = 12'h581;
20'b00000111000000110101 : ColourData = 12'h360;
20'b00000111010000110101 : ColourData = 12'h360;
20'b00000111100000110101 : ColourData = 12'h360;
20'b00000111110000110101 : ColourData = 12'h360;
20'b00001000000000110101 : ColourData = 12'h581;
20'b00001000010000110101 : ColourData = 12'h5A1;
20'b00001000100000110101 : ColourData = 12'h5A1;
20'b00001000110000110101 : ColourData = 12'h5A1;
20'b00001001000000110101 : ColourData = 12'h5A1;
20'b00001001010000110101 : ColourData = 12'h5A1;
20'b00001001100000110101 : ColourData = 12'h5A1;
20'b00001001110000110101 : ColourData = 12'h5A1;
20'b00001010000000110101 : ColourData = 12'h5A1;
20'b00001010010000110101 : ColourData = 12'h5A1;
20'b00001010100000110101 : ColourData = 12'h5A1;
20'b00001010110000110101 : ColourData = 12'h5A1;
20'b00001011000000110101 : ColourData = 12'h5A1;
20'b00001011010000110101 : ColourData = 12'h5A1;
20'b00001011100000110101 : ColourData = 12'h5A1;
20'b00001011110000110101 : ColourData = 12'h6A1;
20'b00001100000000110101 : ColourData = 12'h481;
20'b00001100010000110101 : ColourData = 12'h360;
20'b00001100100000110101 : ColourData = 12'h360;
20'b00001100110000110101 : ColourData = 12'h360;
20'b00001101000000110101 : ColourData = 12'h360;
20'b00001101010000110101 : ColourData = 12'h000;
20'b00001101100000110101 : ColourData = 12'h000;
20'b00001101110000110101 : ColourData = 12'h000;
20'b00001110000000110101 : ColourData = 12'h000;
20'b00001110010000110101 : ColourData = 12'h000;
20'b00001110100000110101 : ColourData = 12'h000;
20'b00001110110000110101 : ColourData = 12'h000;
20'b00000000000000110110 : ColourData = 12'h000;
20'b00000000010000110110 : ColourData = 12'h000;
20'b00000000100000110110 : ColourData = 12'h000;
20'b00000000110000110110 : ColourData = 12'h000;
20'b00000001000000110110 : ColourData = 12'h000;
20'b00000001010000110110 : ColourData = 12'h000;
20'b00000001100000110110 : ColourData = 12'h010;
20'b00000001110000110110 : ColourData = 12'h360;
20'b00000010000000110110 : ColourData = 12'h360;
20'b00000010010000110110 : ColourData = 12'h360;
20'b00000010100000110110 : ColourData = 12'h360;
20'b00000010110000110110 : ColourData = 12'h471;
20'b00000011000000110110 : ColourData = 12'h591;
20'b00000011010000110110 : ColourData = 12'h591;
20'b00000011100000110110 : ColourData = 12'h5A1;
20'b00000011110000110110 : ColourData = 12'h5A1;
20'b00000100000000110110 : ColourData = 12'h5A1;
20'b00000100010000110110 : ColourData = 12'h5A1;
20'b00000100100000110110 : ColourData = 12'h5A1;
20'b00000100110000110110 : ColourData = 12'h5A1;
20'b00000101000000110110 : ColourData = 12'h5A1;
20'b00000101010000110110 : ColourData = 12'h5A1;
20'b00000101100000110110 : ColourData = 12'h5A1;
20'b00000101110000110110 : ColourData = 12'h5A1;
20'b00000110000000110110 : ColourData = 12'h5A1;
20'b00000110010000110110 : ColourData = 12'h5A1;
20'b00000110100000110110 : ColourData = 12'h5A1;
20'b00000110110000110110 : ColourData = 12'h581;
20'b00000111000000110110 : ColourData = 12'h360;
20'b00000111010000110110 : ColourData = 12'h360;
20'b00000111100000110110 : ColourData = 12'h360;
20'b00000111110000110110 : ColourData = 12'h360;
20'b00001000000000110110 : ColourData = 12'h581;
20'b00001000010000110110 : ColourData = 12'h5A1;
20'b00001000100000110110 : ColourData = 12'h5A1;
20'b00001000110000110110 : ColourData = 12'h5A1;
20'b00001001000000110110 : ColourData = 12'h5A1;
20'b00001001010000110110 : ColourData = 12'h5A1;
20'b00001001100000110110 : ColourData = 12'h5A1;
20'b00001001110000110110 : ColourData = 12'h5A1;
20'b00001010000000110110 : ColourData = 12'h5A1;
20'b00001010010000110110 : ColourData = 12'h5A1;
20'b00001010100000110110 : ColourData = 12'h5A1;
20'b00001010110000110110 : ColourData = 12'h5A1;
20'b00001011000000110110 : ColourData = 12'h5A1;
20'b00001011010000110110 : ColourData = 12'h5A1;
20'b00001011100000110110 : ColourData = 12'h591;
20'b00001011110000110110 : ColourData = 12'h591;
20'b00001100000000110110 : ColourData = 12'h471;
20'b00001100010000110110 : ColourData = 12'h360;
20'b00001100100000110110 : ColourData = 12'h360;
20'b00001100110000110110 : ColourData = 12'h360;
20'b00001101000000110110 : ColourData = 12'h360;
20'b00001101010000110110 : ColourData = 12'h010;
20'b00001101100000110110 : ColourData = 12'h000;
20'b00001101110000110110 : ColourData = 12'h000;
20'b00001110000000110110 : ColourData = 12'h000;
20'b00001110010000110110 : ColourData = 12'h000;
20'b00001110100000110110 : ColourData = 12'h000;
20'b00001110110000110110 : ColourData = 12'h000;
20'b00000000000000110111 : ColourData = 12'h333;
20'b00000000010000110111 : ColourData = 12'h333;
20'b00000000100000110111 : ColourData = 12'h333;
20'b00000000110000110111 : ColourData = 12'h333;
20'b00000001000000110111 : ColourData = 12'h333;
20'b00000001010000110111 : ColourData = 12'h333;
20'b00000001100000110111 : ColourData = 12'h333;
20'b00000001110000110111 : ColourData = 12'h360;
20'b00000010000000110111 : ColourData = 12'h360;
20'b00000010010000110111 : ColourData = 12'h360;
20'b00000010100000110111 : ColourData = 12'h360;
20'b00000010110000110111 : ColourData = 12'h360;
20'b00000011000000110111 : ColourData = 12'h350;
20'b00000011010000110111 : ColourData = 12'h360;
20'b00000011100000110111 : ColourData = 12'h5A1;
20'b00000011110000110111 : ColourData = 12'h5A1;
20'b00000100000000110111 : ColourData = 12'h5A1;
20'b00000100010000110111 : ColourData = 12'h5A1;
20'b00000100100000110111 : ColourData = 12'h5A1;
20'b00000100110000110111 : ColourData = 12'h5A1;
20'b00000101000000110111 : ColourData = 12'h5A1;
20'b00000101010000110111 : ColourData = 12'h5A1;
20'b00000101100000110111 : ColourData = 12'h5A1;
20'b00000101110000110111 : ColourData = 12'h5A1;
20'b00000110000000110111 : ColourData = 12'h5A1;
20'b00000110010000110111 : ColourData = 12'h5A1;
20'b00000110100000110111 : ColourData = 12'h6A1;
20'b00000110110000110111 : ColourData = 12'h591;
20'b00000111000000110111 : ColourData = 12'h360;
20'b00000111010000110111 : ColourData = 12'h360;
20'b00000111100000110111 : ColourData = 12'h360;
20'b00000111110000110111 : ColourData = 12'h360;
20'b00001000000000110111 : ColourData = 12'h591;
20'b00001000010000110111 : ColourData = 12'h6A1;
20'b00001000100000110111 : ColourData = 12'h5A1;
20'b00001000110000110111 : ColourData = 12'h5A1;
20'b00001001000000110111 : ColourData = 12'h5A1;
20'b00001001010000110111 : ColourData = 12'h5A1;
20'b00001001100000110111 : ColourData = 12'h5A1;
20'b00001001110000110111 : ColourData = 12'h5A1;
20'b00001010000000110111 : ColourData = 12'h5A1;
20'b00001010010000110111 : ColourData = 12'h5A1;
20'b00001010100000110111 : ColourData = 12'h5A1;
20'b00001010110000110111 : ColourData = 12'h5A1;
20'b00001011000000110111 : ColourData = 12'h5A1;
20'b00001011010000110111 : ColourData = 12'h5A1;
20'b00001011100000110111 : ColourData = 12'h360;
20'b00001011110000110111 : ColourData = 12'h350;
20'b00001100000000110111 : ColourData = 12'h360;
20'b00001100010000110111 : ColourData = 12'h360;
20'b00001100100000110111 : ColourData = 12'h360;
20'b00001100110000110111 : ColourData = 12'h360;
20'b00001101000000110111 : ColourData = 12'h360;
20'b00001101010000110111 : ColourData = 12'h333;
20'b00001101100000110111 : ColourData = 12'h333;
20'b00001101110000110111 : ColourData = 12'h333;
20'b00001110000000110111 : ColourData = 12'h333;
20'b00001110010000110111 : ColourData = 12'h333;
20'b00001110100000110111 : ColourData = 12'h333;
20'b00001110110000110111 : ColourData = 12'h333;
20'b00000000000000111000 : ColourData = 12'hAAA;
20'b00000000010000111000 : ColourData = 12'hAAA;
20'b00000000100000111000 : ColourData = 12'hAAA;
20'b00000000110000111000 : ColourData = 12'hAAA;
20'b00000001000000111000 : ColourData = 12'hAAA;
20'b00000001010000111000 : ColourData = 12'hAAA;
20'b00000001100000111000 : ColourData = 12'h999;
20'b00000001110000111000 : ColourData = 12'h360;
20'b00000010000000111000 : ColourData = 12'h360;
20'b00000010010000111000 : ColourData = 12'h360;
20'b00000010100000111000 : ColourData = 12'h360;
20'b00000010110000111000 : ColourData = 12'h360;
20'b00000011000000111000 : ColourData = 12'h360;
20'b00000011010000111000 : ColourData = 12'h360;
20'b00000011100000111000 : ColourData = 12'h481;
20'b00000011110000111000 : ColourData = 12'h481;
20'b00000100000000111000 : ColourData = 12'h481;
20'b00000100010000111000 : ColourData = 12'h481;
20'b00000100100000111000 : ColourData = 12'h481;
20'b00000100110000111000 : ColourData = 12'h481;
20'b00000101000000111000 : ColourData = 12'h481;
20'b00000101010000111000 : ColourData = 12'h481;
20'b00000101100000111000 : ColourData = 12'h481;
20'b00000101110000111000 : ColourData = 12'h481;
20'b00000110000000111000 : ColourData = 12'h481;
20'b00000110010000111000 : ColourData = 12'h481;
20'b00000110100000111000 : ColourData = 12'h481;
20'b00000110110000111000 : ColourData = 12'h471;
20'b00000111000000111000 : ColourData = 12'h360;
20'b00000111010000111000 : ColourData = 12'h360;
20'b00000111100000111000 : ColourData = 12'h360;
20'b00000111110000111000 : ColourData = 12'h360;
20'b00001000000000111000 : ColourData = 12'h471;
20'b00001000010000111000 : ColourData = 12'h481;
20'b00001000100000111000 : ColourData = 12'h481;
20'b00001000110000111000 : ColourData = 12'h481;
20'b00001001000000111000 : ColourData = 12'h481;
20'b00001001010000111000 : ColourData = 12'h481;
20'b00001001100000111000 : ColourData = 12'h481;
20'b00001001110000111000 : ColourData = 12'h481;
20'b00001010000000111000 : ColourData = 12'h481;
20'b00001010010000111000 : ColourData = 12'h481;
20'b00001010100000111000 : ColourData = 12'h481;
20'b00001010110000111000 : ColourData = 12'h481;
20'b00001011000000111000 : ColourData = 12'h481;
20'b00001011010000111000 : ColourData = 12'h481;
20'b00001011100000111000 : ColourData = 12'h360;
20'b00001011110000111000 : ColourData = 12'h360;
20'b00001100000000111000 : ColourData = 12'h360;
20'b00001100010000111000 : ColourData = 12'h360;
20'b00001100100000111000 : ColourData = 12'h360;
20'b00001100110000111000 : ColourData = 12'h360;
20'b00001101000000111000 : ColourData = 12'h360;
20'b00001101010000111000 : ColourData = 12'h999;
20'b00001101100000111000 : ColourData = 12'hAAA;
20'b00001101110000111000 : ColourData = 12'hAAA;
20'b00001110000000111000 : ColourData = 12'hAAA;
20'b00001110010000111000 : ColourData = 12'hAAA;
20'b00001110100000111000 : ColourData = 12'hAAA;
20'b00001110110000111000 : ColourData = 12'hAAA;
20'b00000000000000111001 : ColourData = 12'hFFF;
20'b00000000010000111001 : ColourData = 12'hFFF;
20'b00000000100000111001 : ColourData = 12'hFFF;
20'b00000000110000111001 : ColourData = 12'hFFF;
20'b00000001000000111001 : ColourData = 12'hFFF;
20'b00000001010000111001 : ColourData = 12'hFFF;
20'b00000001100000111001 : ColourData = 12'hEEE;
20'b00000001110000111001 : ColourData = 12'h250;
20'b00000010000000111001 : ColourData = 12'h250;
20'b00000010010000111001 : ColourData = 12'h360;
20'b00000010100000111001 : ColourData = 12'h360;
20'b00000010110000111001 : ColourData = 12'h360;
20'b00000011000000111001 : ColourData = 12'h360;
20'b00000011010000111001 : ColourData = 12'h360;
20'b00000011100000111001 : ColourData = 12'h360;
20'b00000011110000111001 : ColourData = 12'h360;
20'b00000100000000111001 : ColourData = 12'h360;
20'b00000100010000111001 : ColourData = 12'h360;
20'b00000100100000111001 : ColourData = 12'h360;
20'b00000100110000111001 : ColourData = 12'h360;
20'b00000101000000111001 : ColourData = 12'h360;
20'b00000101010000111001 : ColourData = 12'h360;
20'b00000101100000111001 : ColourData = 12'h360;
20'b00000101110000111001 : ColourData = 12'h360;
20'b00000110000000111001 : ColourData = 12'h360;
20'b00000110010000111001 : ColourData = 12'h360;
20'b00000110100000111001 : ColourData = 12'h360;
20'b00000110110000111001 : ColourData = 12'h360;
20'b00000111000000111001 : ColourData = 12'h360;
20'b00000111010000111001 : ColourData = 12'h360;
20'b00000111100000111001 : ColourData = 12'h360;
20'b00000111110000111001 : ColourData = 12'h360;
20'b00001000000000111001 : ColourData = 12'h360;
20'b00001000010000111001 : ColourData = 12'h360;
20'b00001000100000111001 : ColourData = 12'h360;
20'b00001000110000111001 : ColourData = 12'h360;
20'b00001001000000111001 : ColourData = 12'h360;
20'b00001001010000111001 : ColourData = 12'h360;
20'b00001001100000111001 : ColourData = 12'h360;
20'b00001001110000111001 : ColourData = 12'h360;
20'b00001010000000111001 : ColourData = 12'h360;
20'b00001010010000111001 : ColourData = 12'h360;
20'b00001010100000111001 : ColourData = 12'h360;
20'b00001010110000111001 : ColourData = 12'h360;
20'b00001011000000111001 : ColourData = 12'h360;
20'b00001011010000111001 : ColourData = 12'h360;
20'b00001011100000111001 : ColourData = 12'h360;
20'b00001011110000111001 : ColourData = 12'h360;
20'b00001100000000111001 : ColourData = 12'h360;
20'b00001100010000111001 : ColourData = 12'h360;
20'b00001100100000111001 : ColourData = 12'h360;
20'b00001100110000111001 : ColourData = 12'h250;
20'b00001101000000111001 : ColourData = 12'h250;
20'b00001101010000111001 : ColourData = 12'hEEE;
20'b00001101100000111001 : ColourData = 12'hFFF;
20'b00001101110000111001 : ColourData = 12'hFFF;
20'b00001110000000111001 : ColourData = 12'hFFF;
20'b00001110010000111001 : ColourData = 12'hFFF;
20'b00001110100000111001 : ColourData = 12'hFFF;
20'b00001110110000111001 : ColourData = 12'hFFF;
20'b00000000000000111010 : ColourData = 12'hFFF;
20'b00000000010000111010 : ColourData = 12'hFFF;
20'b00000000100000111010 : ColourData = 12'hFFF;
20'b00000000110000111010 : ColourData = 12'hFFF;
20'b00000001000000111010 : ColourData = 12'hFFF;
20'b00000001010000111010 : ColourData = 12'hFFF;
20'b00000001100000111010 : ColourData = 12'hFFF;
20'b00000001110000111010 : ColourData = 12'hDDC;
20'b00000010000000111010 : ColourData = 12'hDDD;
20'b00000010010000111010 : ColourData = 12'h573;
20'b00000010100000111010 : ColourData = 12'h360;
20'b00000010110000111010 : ColourData = 12'h360;
20'b00000011000000111010 : ColourData = 12'h360;
20'b00000011010000111010 : ColourData = 12'h360;
20'b00000011100000111010 : ColourData = 12'h360;
20'b00000011110000111010 : ColourData = 12'h360;
20'b00000100000000111010 : ColourData = 12'h360;
20'b00000100010000111010 : ColourData = 12'h360;
20'b00000100100000111010 : ColourData = 12'h360;
20'b00000100110000111010 : ColourData = 12'h360;
20'b00000101000000111010 : ColourData = 12'h360;
20'b00000101010000111010 : ColourData = 12'h360;
20'b00000101100000111010 : ColourData = 12'h360;
20'b00000101110000111010 : ColourData = 12'h360;
20'b00000110000000111010 : ColourData = 12'h360;
20'b00000110010000111010 : ColourData = 12'h360;
20'b00000110100000111010 : ColourData = 12'h360;
20'b00000110110000111010 : ColourData = 12'h360;
20'b00000111000000111010 : ColourData = 12'h360;
20'b00000111010000111010 : ColourData = 12'h360;
20'b00000111100000111010 : ColourData = 12'h360;
20'b00000111110000111010 : ColourData = 12'h360;
20'b00001000000000111010 : ColourData = 12'h360;
20'b00001000010000111010 : ColourData = 12'h360;
20'b00001000100000111010 : ColourData = 12'h360;
20'b00001000110000111010 : ColourData = 12'h360;
20'b00001001000000111010 : ColourData = 12'h360;
20'b00001001010000111010 : ColourData = 12'h360;
20'b00001001100000111010 : ColourData = 12'h360;
20'b00001001110000111010 : ColourData = 12'h360;
20'b00001010000000111010 : ColourData = 12'h360;
20'b00001010010000111010 : ColourData = 12'h360;
20'b00001010100000111010 : ColourData = 12'h360;
20'b00001010110000111010 : ColourData = 12'h360;
20'b00001011000000111010 : ColourData = 12'h360;
20'b00001011010000111010 : ColourData = 12'h360;
20'b00001011100000111010 : ColourData = 12'h360;
20'b00001011110000111010 : ColourData = 12'h360;
20'b00001100000000111010 : ColourData = 12'h360;
20'b00001100010000111010 : ColourData = 12'h360;
20'b00001100100000111010 : ColourData = 12'h573;
20'b00001100110000111010 : ColourData = 12'hDDD;
20'b00001101000000111010 : ColourData = 12'hDDC;
20'b00001101010000111010 : ColourData = 12'hFFF;
20'b00001101100000111010 : ColourData = 12'hFFF;
20'b00001101110000111010 : ColourData = 12'hFFF;
20'b00001110000000111010 : ColourData = 12'hFFF;
20'b00001110010000111010 : ColourData = 12'hFFF;
20'b00001110100000111010 : ColourData = 12'hFFF;
20'b00001110110000111010 : ColourData = 12'hFFF;
20'b00000000000000111011 : ColourData = 12'hFFF;
20'b00000000010000111011 : ColourData = 12'hFFF;
20'b00000000100000111011 : ColourData = 12'hFFF;
20'b00000000110000111011 : ColourData = 12'hFFF;
20'b00000001000000111011 : ColourData = 12'hFFF;
20'b00000001010000111011 : ColourData = 12'hFFF;
20'b00000001100000111011 : ColourData = 12'hFFF;
20'b00000001110000111011 : ColourData = 12'hFFF;
20'b00000010000000111011 : ColourData = 12'hFFF;
20'b00000010010000111011 : ColourData = 12'h684;
20'b00000010100000111011 : ColourData = 12'h350;
20'b00000010110000111011 : ColourData = 12'h360;
20'b00000011000000111011 : ColourData = 12'h360;
20'b00000011010000111011 : ColourData = 12'h360;
20'b00000011100000111011 : ColourData = 12'h360;
20'b00000011110000111011 : ColourData = 12'h360;
20'b00000100000000111011 : ColourData = 12'h360;
20'b00000100010000111011 : ColourData = 12'h360;
20'b00000100100000111011 : ColourData = 12'h360;
20'b00000100110000111011 : ColourData = 12'h360;
20'b00000101000000111011 : ColourData = 12'h360;
20'b00000101010000111011 : ColourData = 12'h360;
20'b00000101100000111011 : ColourData = 12'h360;
20'b00000101110000111011 : ColourData = 12'h360;
20'b00000110000000111011 : ColourData = 12'h360;
20'b00000110010000111011 : ColourData = 12'h360;
20'b00000110100000111011 : ColourData = 12'h360;
20'b00000110110000111011 : ColourData = 12'h360;
20'b00000111000000111011 : ColourData = 12'h360;
20'b00000111010000111011 : ColourData = 12'h360;
20'b00000111100000111011 : ColourData = 12'h360;
20'b00000111110000111011 : ColourData = 12'h360;
20'b00001000000000111011 : ColourData = 12'h360;
20'b00001000010000111011 : ColourData = 12'h360;
20'b00001000100000111011 : ColourData = 12'h360;
20'b00001000110000111011 : ColourData = 12'h360;
20'b00001001000000111011 : ColourData = 12'h360;
20'b00001001010000111011 : ColourData = 12'h360;
20'b00001001100000111011 : ColourData = 12'h360;
20'b00001001110000111011 : ColourData = 12'h360;
20'b00001010000000111011 : ColourData = 12'h360;
20'b00001010010000111011 : ColourData = 12'h360;
20'b00001010100000111011 : ColourData = 12'h360;
20'b00001010110000111011 : ColourData = 12'h360;
20'b00001011000000111011 : ColourData = 12'h360;
20'b00001011010000111011 : ColourData = 12'h360;
20'b00001011100000111011 : ColourData = 12'h360;
20'b00001011110000111011 : ColourData = 12'h360;
20'b00001100000000111011 : ColourData = 12'h360;
20'b00001100010000111011 : ColourData = 12'h350;
20'b00001100100000111011 : ColourData = 12'h684;
20'b00001100110000111011 : ColourData = 12'hFFF;
20'b00001101000000111011 : ColourData = 12'hFFF;
20'b00001101010000111011 : ColourData = 12'hFFF;
20'b00001101100000111011 : ColourData = 12'hFFF;
20'b00001101110000111011 : ColourData = 12'hFFF;
20'b00001110000000111011 : ColourData = 12'hFFF;
20'b00001110010000111011 : ColourData = 12'hFFF;
20'b00001110100000111011 : ColourData = 12'hFFF;
20'b00001110110000111011 : ColourData = 12'hFFF;


default: ColourData = 12'h000;

endcase
end

endmodule
