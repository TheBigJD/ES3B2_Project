module Bottle(
input Master_Clock_In,
input [9 : 0] xInput,
input [9 : 0] yInput,
output reg [11:0] ColourData = 12'h000
//output reg [3:0] Red_Out, Green_Out, Blue_Out = 4'h0
);

(* rom_style = "block" *)

//reg [11:0] ColourData;
reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

//reg [11:0] ColourData = 12'h000;

always @(posedge Master_Clock_In)
begin


a = xInput % 32;
b = yInput % 160;

Inputs = {a, b};

	//if ((x < 640) & (y < 480)) begin
    case(Inputs)

20'b00000000000000000000:ColourData=12'h964;
20'b00000000010000000000:ColourData=12'hB65;
20'b00000000100000000000:ColourData=12'hC77;
20'b00000000110000000000:ColourData=12'hC76;
20'b00000001000000000000:ColourData=12'hC76;
20'b00000001010000000000:ColourData=12'hC76;
20'b00000001100000000000:ColourData=12'hC77;
20'b00000001110000000000:ColourData=12'hB66;
20'b00000010000000000000:ColourData=12'h211;
20'b00000010010000000000:ColourData=12'hB66;
20'b00000010100000000000:ColourData=12'hC77;
20'b00000010110000000000:ColourData=12'hC76;
20'b00000011000000000000:ColourData=12'hC76;
20'b00000011010000000000:ColourData=12'hC77;
20'b00000011100000000000:ColourData=12'hB65;
20'b00000011110000000000:ColourData=12'h773;
20'b00000100000000000000:ColourData=12'h0F0;
20'b00000100010000000000:ColourData=12'h0F0;
20'b00000100100000000000:ColourData=12'h0F0;
20'b00000100110000000000:ColourData=12'h0F0;
20'b00000101000000000000:ColourData=12'h0F0;
20'b00000101010000000000:ColourData=12'h5B0;
20'b00000101100000000000:ColourData=12'hD50;
20'b00000101110000000000:ColourData=12'hD40;
20'b00000110000000000000:ColourData=12'hE40;
20'b00000110010000000000:ColourData=12'hA70;
20'b00000110100000000000:ColourData=12'h1E0;
20'b00000110110000000000:ColourData=12'h0F0;
20'b00000111000000000000:ColourData=12'h0F0;
20'b00000111010000000000:ColourData=12'h0F0;
20'b00000111100000000000:ColourData=12'h0F0;
20'b00000111110000000000:ColourData=12'h6F6;
20'b00000000000000000001:ColourData=12'hD88;
20'b00000000010000000001:ColourData=12'h842;
20'b00000000100000000001:ColourData=12'h731;
20'b00000000110000000001:ColourData=12'h731;
20'b00000001000000000001:ColourData=12'h731;
20'b00000001010000000001:ColourData=12'h731;
20'b00000001100000000001:ColourData=12'h741;
20'b00000001110000000001:ColourData=12'h730;
20'b00000010000000000001:ColourData=12'h100;
20'b00000010010000000001:ColourData=12'hA66;
20'b00000010100000000001:ColourData=12'h842;
20'b00000010110000000001:ColourData=12'h731;
20'b00000011000000000001:ColourData=12'h731;
20'b00000011010000000001:ColourData=12'h741;
20'b00000011100000000001:ColourData=12'h620;
20'b00000011110000000001:ColourData=12'h342;
20'b00000100000000000001:ColourData=12'h0F0;
20'b00000100010000000001:ColourData=12'h0F0;
20'b00000100100000000001:ColourData=12'h0F0;
20'b00000100110000000001:ColourData=12'h0F0;
20'b00000101000000000001:ColourData=12'h5B0;
20'b00000101010000000001:ColourData=12'hD50;
20'b00000101100000000001:ColourData=12'hD40;
20'b00000101110000000001:ColourData=12'hD50;
20'b00000110000000000001:ColourData=12'hD50;
20'b00000110010000000001:ColourData=12'hE40;
20'b00000110100000000001:ColourData=12'hA70;
20'b00000110110000000001:ColourData=12'h1E0;
20'b00000111000000000001:ColourData=12'h0F0;
20'b00000111010000000001:ColourData=12'h0F0;
20'b00000111100000000001:ColourData=12'h0F0;
20'b00000111110000000001:ColourData=12'h6F6;
20'b00000000000000000010:ColourData=12'hD99;
20'b00000000010000000010:ColourData=12'h841;
20'b00000000100000000010:ColourData=12'h730;
20'b00000000110000000010:ColourData=12'h730;
20'b00000001000000000010:ColourData=12'h730;
20'b00000001010000000010:ColourData=12'h730;
20'b00000001100000000010:ColourData=12'h730;
20'b00000001110000000010:ColourData=12'h630;
20'b00000010000000000010:ColourData=12'h100;
20'b00000010010000000010:ColourData=12'hA65;
20'b00000010100000000010:ColourData=12'h841;
20'b00000010110000000010:ColourData=12'h730;
20'b00000011000000000010:ColourData=12'h730;
20'b00000011010000000010:ColourData=12'h730;
20'b00000011100000000010:ColourData=12'h520;
20'b00000011110000000010:ColourData=12'h242;
20'b00000100000000000010:ColourData=12'h0F0;
20'b00000100010000000010:ColourData=12'h0F0;
20'b00000100100000000010:ColourData=12'h0F0;
20'b00000100110000000010:ColourData=12'h5B0;
20'b00000101000000000010:ColourData=12'hD50;
20'b00000101010000000010:ColourData=12'hD40;
20'b00000101100000000010:ColourData=12'hD50;
20'b00000101110000000010:ColourData=12'hD50;
20'b00000110000000000010:ColourData=12'hD50;
20'b00000110010000000010:ColourData=12'hD50;
20'b00000110100000000010:ColourData=12'hE40;
20'b00000110110000000010:ColourData=12'hA70;
20'b00000111000000000010:ColourData=12'h1E0;
20'b00000111010000000010:ColourData=12'h0F0;
20'b00000111100000000010:ColourData=12'h0F0;
20'b00000111110000000010:ColourData=12'h6F6;
20'b00000000000000000011:ColourData=12'hD99;
20'b00000000010000000011:ColourData=12'h841;
20'b00000000100000000011:ColourData=12'h730;
20'b00000000110000000011:ColourData=12'h730;
20'b00000001000000000011:ColourData=12'h730;
20'b00000001010000000011:ColourData=12'h730;
20'b00000001100000000011:ColourData=12'h730;
20'b00000001110000000011:ColourData=12'h630;
20'b00000010000000000011:ColourData=12'h100;
20'b00000010010000000011:ColourData=12'hA66;
20'b00000010100000000011:ColourData=12'h731;
20'b00000010110000000011:ColourData=12'h730;
20'b00000011000000000011:ColourData=12'h730;
20'b00000011010000000011:ColourData=12'h730;
20'b00000011100000000011:ColourData=12'h620;
20'b00000011110000000011:ColourData=12'h242;
20'b00000100000000000011:ColourData=12'h0F0;
20'b00000100010000000011:ColourData=12'h0F0;
20'b00000100100000000011:ColourData=12'h4B0;
20'b00000100110000000011:ColourData=12'hA40;
20'b00000101000000000011:ColourData=12'hB40;
20'b00000101010000000011:ColourData=12'hE50;
20'b00000101100000000011:ColourData=12'hD50;
20'b00000101110000000011:ColourData=12'hD50;
20'b00000110000000000011:ColourData=12'hD50;
20'b00000110010000000011:ColourData=12'hE50;
20'b00000110100000000011:ColourData=12'hC40;
20'b00000110110000000011:ColourData=12'hA30;
20'b00000111000000000011:ColourData=12'h770;
20'b00000111010000000011:ColourData=12'h1E0;
20'b00000111100000000011:ColourData=12'h0F0;
20'b00000111110000000011:ColourData=12'h6F6;
20'b00000000000000000100:ColourData=12'hD99;
20'b00000000010000000100:ColourData=12'h841;
20'b00000000100000000100:ColourData=12'h730;
20'b00000000110000000100:ColourData=12'h730;
20'b00000001000000000100:ColourData=12'h730;
20'b00000001010000000100:ColourData=12'h730;
20'b00000001100000000100:ColourData=12'h730;
20'b00000001110000000100:ColourData=12'h630;
20'b00000010000000000100:ColourData=12'h100;
20'b00000010010000000100:ColourData=12'h955;
20'b00000010100000000100:ColourData=12'h210;
20'b00000010110000000100:ColourData=12'h520;
20'b00000011000000000100:ColourData=12'h630;
20'b00000011010000000100:ColourData=12'h630;
20'b00000011100000000100:ColourData=12'h520;
20'b00000011110000000100:ColourData=12'h342;
20'b00000100000000000100:ColourData=12'h0F0;
20'b00000100010000000100:ColourData=12'h5B0;
20'b00000100100000000100:ColourData=12'hB40;
20'b00000100110000000100:ColourData=12'h421;
20'b00000101000000000100:ColourData=12'h642;
20'b00000101010000000100:ColourData=12'hB40;
20'b00000101100000000100:ColourData=12'hE50;
20'b00000101110000000100:ColourData=12'hE50;
20'b00000110000000000100:ColourData=12'hE50;
20'b00000110010000000100:ColourData=12'hD40;
20'b00000110100000000100:ColourData=12'h841;
20'b00000110110000000100:ColourData=12'h432;
20'b00000111000000000100:ColourData=12'h820;
20'b00000111010000000100:ColourData=12'h980;
20'b00000111100000000100:ColourData=12'h1E0;
20'b00000111110000000100:ColourData=12'h6F6;
20'b00000000000000000101:ColourData=12'hD99;
20'b00000000010000000101:ColourData=12'h841;
20'b00000000100000000101:ColourData=12'h730;
20'b00000000110000000101:ColourData=12'h730;
20'b00000001000000000101:ColourData=12'h730;
20'b00000001010000000101:ColourData=12'h730;
20'b00000001100000000101:ColourData=12'h730;
20'b00000001110000000101:ColourData=12'h630;
20'b00000010000000000101:ColourData=12'h100;
20'b00000010010000000101:ColourData=12'h631;
20'b00000010100000000101:ColourData=12'h100;
20'b00000010110000000101:ColourData=12'h100;
20'b00000011000000000101:ColourData=12'h100;
20'b00000011010000000101:ColourData=12'h100;
20'b00000011100000000101:ColourData=12'h200;
20'b00000011110000000101:ColourData=12'h562;
20'b00000100000000000101:ColourData=12'h2D0;
20'b00000100010000000101:ColourData=12'hD50;
20'b00000100100000000101:ColourData=12'hD40;
20'b00000100110000000101:ColourData=12'hE73;
20'b00000101000000000101:ColourData=12'hB98;
20'b00000101010000000101:ColourData=12'h321;
20'b00000101100000000101:ColourData=12'hA30;
20'b00000101110000000101:ColourData=12'hA40;
20'b00000110000000000101:ColourData=12'hA40;
20'b00000110010000000101:ColourData=12'h720;
20'b00000110100000000101:ColourData=12'h554;
20'b00000110110000000101:ColourData=12'hEA7;
20'b00000111000000000101:ColourData=12'hD40;
20'b00000111010000000101:ColourData=12'hE40;
20'b00000111100000000101:ColourData=12'h790;
20'b00000111110000000101:ColourData=12'h5F6;
20'b00000000000000000110:ColourData=12'hD99;
20'b00000000010000000110:ColourData=12'h841;
20'b00000000100000000110:ColourData=12'h730;
20'b00000000110000000110:ColourData=12'h730;
20'b00000001000000000110:ColourData=12'h730;
20'b00000001010000000110:ColourData=12'h730;
20'b00000001100000000110:ColourData=12'h730;
20'b00000001110000000110:ColourData=12'h630;
20'b00000010000000000110:ColourData=12'h100;
20'b00000010010000000110:ColourData=12'hA55;
20'b00000010100000000110:ColourData=12'hB66;
20'b00000010110000000110:ColourData=12'hB66;
20'b00000011000000000110:ColourData=12'hB66;
20'b00000011010000000110:ColourData=12'hB66;
20'b00000011100000000110:ColourData=12'h945;
20'b00000011110000000110:ColourData=12'h342;
20'b00000100000000000110:ColourData=12'h5B0;
20'b00000100010000000110:ColourData=12'hD50;
20'b00000100100000000110:ColourData=12'hD40;
20'b00000100110000000110:ColourData=12'hE73;
20'b00000101000000000110:ColourData=12'hB98;
20'b00000101010000000110:ColourData=12'h222;
20'b00000101100000000110:ColourData=12'h432;
20'b00000101110000000110:ColourData=12'h421;
20'b00000110000000000110:ColourData=12'h422;
20'b00000110010000000110:ColourData=12'h322;
20'b00000110100000000110:ColourData=12'h554;
20'b00000110110000000110:ColourData=12'hEA7;
20'b00000111000000000110:ColourData=12'hD40;
20'b00000111010000000110:ColourData=12'hE40;
20'b00000111100000000110:ColourData=12'h970;
20'b00000111110000000110:ColourData=12'h7E6;
20'b00000000000000000111:ColourData=12'hD99;
20'b00000000010000000111:ColourData=12'h841;
20'b00000000100000000111:ColourData=12'h730;
20'b00000000110000000111:ColourData=12'h730;
20'b00000001000000000111:ColourData=12'h730;
20'b00000001010000000111:ColourData=12'h730;
20'b00000001100000000111:ColourData=12'h730;
20'b00000001110000000111:ColourData=12'h630;
20'b00000010000000000111:ColourData=12'h100;
20'b00000010010000000111:ColourData=12'hA66;
20'b00000010100000000111:ColourData=12'h842;
20'b00000010110000000111:ColourData=12'h741;
20'b00000011000000000111:ColourData=12'h741;
20'b00000011010000000111:ColourData=12'h841;
20'b00000011100000000111:ColourData=12'h630;
20'b00000011110000000111:ColourData=12'h432;
20'b00000100000000000111:ColourData=12'hD51;
20'b00000100010000000111:ColourData=12'hD40;
20'b00000100100000000111:ColourData=12'hD40;
20'b00000100110000000111:ColourData=12'hE73;
20'b00000101000000000111:ColourData=12'hCA9;
20'b00000101010000000111:ColourData=12'h766;
20'b00000101100000000111:ColourData=12'hEA8;
20'b00000101110000000111:ColourData=12'hD40;
20'b00000110000000000111:ColourData=12'hE73;
20'b00000110010000000111:ColourData=12'hB98;
20'b00000110100000000111:ColourData=12'h776;
20'b00000110110000000111:ColourData=12'hEA7;
20'b00000111000000000111:ColourData=12'hD40;
20'b00000111010000000111:ColourData=12'hD50;
20'b00000111100000000111:ColourData=12'hD40;
20'b00000111110000000111:ColourData=12'hE96;
20'b00000000000000001000:ColourData=12'hD99;
20'b00000000010000001000:ColourData=12'h841;
20'b00000000100000001000:ColourData=12'h730;
20'b00000000110000001000:ColourData=12'h730;
20'b00000001000000001000:ColourData=12'h730;
20'b00000001010000001000:ColourData=12'h730;
20'b00000001100000001000:ColourData=12'h730;
20'b00000001110000001000:ColourData=12'h630;
20'b00000010000000001000:ColourData=12'h100;
20'b00000010010000001000:ColourData=12'hA66;
20'b00000010100000001000:ColourData=12'h841;
20'b00000010110000001000:ColourData=12'h730;
20'b00000011000000001000:ColourData=12'h730;
20'b00000011010000001000:ColourData=12'h730;
20'b00000011100000001000:ColourData=12'h520;
20'b00000011110000001000:ColourData=12'h432;
20'b00000100000000001000:ColourData=12'hE51;
20'b00000100010000001000:ColourData=12'hD40;
20'b00000100100000001000:ColourData=12'hD40;
20'b00000100110000001000:ColourData=12'hD62;
20'b00000101000000001000:ColourData=12'hEA8;
20'b00000101010000001000:ColourData=12'hEA8;
20'b00000101100000001000:ColourData=12'hE96;
20'b00000101110000001000:ColourData=12'hD40;
20'b00000110000000001000:ColourData=12'hE62;
20'b00000110010000001000:ColourData=12'hEA8;
20'b00000110100000001000:ColourData=12'hEB8;
20'b00000110110000001000:ColourData=12'hE85;
20'b00000111000000001000:ColourData=12'hD40;
20'b00000111010000001000:ColourData=12'hD50;
20'b00000111100000001000:ColourData=12'hD40;
20'b00000111110000001000:ColourData=12'hE96;
20'b00000000000000001001:ColourData=12'hC88;
20'b00000000010000001001:ColourData=12'h731;
20'b00000000100000001001:ColourData=12'h730;
20'b00000000110000001001:ColourData=12'h730;
20'b00000001000000001001:ColourData=12'h730;
20'b00000001010000001001:ColourData=12'h730;
20'b00000001100000001001:ColourData=12'h730;
20'b00000001110000001001:ColourData=12'h630;
20'b00000010000000001001:ColourData=12'h210;
20'b00000010010000001001:ColourData=12'hA55;
20'b00000010100000001001:ColourData=12'h841;
20'b00000010110000001001:ColourData=12'h730;
20'b00000011000000001001:ColourData=12'h730;
20'b00000011010000001001:ColourData=12'h730;
20'b00000011100000001001:ColourData=12'h520;
20'b00000011110000001001:ColourData=12'h332;
20'b00000100000000001001:ColourData=12'hB71;
20'b00000100010000001001:ColourData=12'hE40;
20'b00000100100000001001:ColourData=12'hE40;
20'b00000100110000001001:ColourData=12'hE40;
20'b00000101000000001001:ColourData=12'hD51;
20'b00000101010000001001:ColourData=12'hE63;
20'b00000101100000001001:ColourData=12'hE62;
20'b00000101110000001001:ColourData=12'hE62;
20'b00000110000000001001:ColourData=12'hD62;
20'b00000110010000001001:ColourData=12'hE63;
20'b00000110100000001001:ColourData=12'hD62;
20'b00000110110000001001:ColourData=12'hD40;
20'b00000111000000001001:ColourData=12'hE40;
20'b00000111010000001001:ColourData=12'hE40;
20'b00000111100000001001:ColourData=12'hC50;
20'b00000111110000001001:ColourData=12'hCA6;
20'b00000000000000001010:ColourData=12'h444;
20'b00000000010000001010:ColourData=12'h100;
20'b00000000100000001010:ColourData=12'h520;
20'b00000000110000001010:ColourData=12'h630;
20'b00000001000000001010:ColourData=12'h730;
20'b00000001010000001010:ColourData=12'h730;
20'b00000001100000001010:ColourData=12'h630;
20'b00000001110000001010:ColourData=12'h100;
20'b00000010000000001010:ColourData=12'h955;
20'b00000010010000001010:ColourData=12'h841;
20'b00000010100000001010:ColourData=12'h730;
20'b00000010110000001010:ColourData=12'h730;
20'b00000011000000001010:ColourData=12'h730;
20'b00000011010000001010:ColourData=12'h730;
20'b00000011100000001010:ColourData=12'h620;
20'b00000011110000001010:ColourData=12'h242;
20'b00000100000000001010:ColourData=12'h2E0;
20'b00000100010000001010:ColourData=12'hA70;
20'b00000100100000001010:ColourData=12'hA70;
20'b00000100110000001010:ColourData=12'hB70;
20'b00000101000000001010:ColourData=12'hE84;
20'b00000101010000001010:ColourData=12'hECA;
20'b00000101100000001010:ColourData=12'hECA;
20'b00000101110000001010:ColourData=12'hECA;
20'b00000110000000001010:ColourData=12'hECA;
20'b00000110010000001010:ColourData=12'hECA;
20'b00000110100000001010:ColourData=12'hEA8;
20'b00000110110000001010:ColourData=12'hC61;
20'b00000111000000001010:ColourData=12'hA70;
20'b00000111010000001010:ColourData=12'hA70;
20'b00000111100000001010:ColourData=12'h5A0;
20'b00000111110000001010:ColourData=12'h6F6;
20'b00000000000000001011:ColourData=12'hC88;
20'b00000000010000001011:ColourData=12'hA55;
20'b00000000100000001011:ColourData=12'h311;
20'b00000000110000001011:ColourData=12'h100;
20'b00000001000000001011:ColourData=12'h520;
20'b00000001010000001011:ColourData=12'h630;
20'b00000001100000001011:ColourData=12'h630;
20'b00000001110000001011:ColourData=12'h210;
20'b00000010000000001011:ColourData=12'hA55;
20'b00000010010000001011:ColourData=12'h841;
20'b00000010100000001011:ColourData=12'h730;
20'b00000010110000001011:ColourData=12'h730;
20'b00000011000000001011:ColourData=12'h730;
20'b00000011010000001011:ColourData=12'h730;
20'b00000011100000001011:ColourData=12'h620;
20'b00000011110000001011:ColourData=12'h242;
20'b00000100000000001011:ColourData=12'h0F0;
20'b00000100010000001011:ColourData=12'h0F0;
20'b00000100100000001011:ColourData=12'h0C0;
20'b00000100110000001011:ColourData=12'h3C2;
20'b00000101000000001011:ColourData=12'hFDA;
20'b00000101010000001011:ColourData=12'hFDB;
20'b00000101100000001011:ColourData=12'hECA;
20'b00000101110000001011:ColourData=12'hECA;
20'b00000110000000001011:ColourData=12'hECA;
20'b00000110010000001011:ColourData=12'hECA;
20'b00000110100000001011:ColourData=12'hFCB;
20'b00000110110000001011:ColourData=12'h9D7;
20'b00000111000000001011:ColourData=12'h0F0;
20'b00000111010000001011:ColourData=12'h0F0;
20'b00000111100000001011:ColourData=12'h0F0;
20'b00000111110000001011:ColourData=12'h6F6;
20'b00000000000000001100:ColourData=12'hD99;
20'b00000000010000001100:ColourData=12'h942;
20'b00000000100000001100:ColourData=12'hA54;
20'b00000000110000001100:ColourData=12'hA66;
20'b00000001000000001100:ColourData=12'h311;
20'b00000001010000001100:ColourData=12'h100;
20'b00000001100000001100:ColourData=12'h100;
20'b00000001110000001100:ColourData=12'h955;
20'b00000010000000001100:ColourData=12'h842;
20'b00000010010000001100:ColourData=12'h730;
20'b00000010100000001100:ColourData=12'h730;
20'b00000010110000001100:ColourData=12'h730;
20'b00000011000000001100:ColourData=12'h730;
20'b00000011010000001100:ColourData=12'h730;
20'b00000011100000001100:ColourData=12'h620;
20'b00000011110000001100:ColourData=12'h242;
20'b00000100000000001100:ColourData=12'h0F0;
20'b00000100010000001100:ColourData=12'h0A0;
20'b00000100100000001100:ColourData=12'h111;
20'b00000100110000001100:ColourData=12'h333;
20'b00000101000000001100:ColourData=12'hBA8;
20'b00000101010000001100:ColourData=12'hCA9;
20'b00000101100000001100:ColourData=12'hFDA;
20'b00000101110000001100:ColourData=12'hECA;
20'b00000110000000001100:ColourData=12'hECA;
20'b00000110010000001100:ColourData=12'hFCA;
20'b00000110100000001100:ColourData=12'hECA;
20'b00000110110000001100:ColourData=12'h7A5;
20'b00000111000000001100:ColourData=12'h0D0;
20'b00000111010000001100:ColourData=12'h0F0;
20'b00000111100000001100:ColourData=12'h0F0;
20'b00000111110000001100:ColourData=12'h6F6;
20'b00000000000000001101:ColourData=12'hD99;
20'b00000000010000001101:ColourData=12'h841;
20'b00000000100000001101:ColourData=12'h730;
20'b00000000110000001101:ColourData=12'h841;
20'b00000001000000001101:ColourData=12'hA55;
20'b00000001010000001101:ColourData=12'hA55;
20'b00000001100000001101:ColourData=12'h101;
20'b00000001110000001101:ColourData=12'hA55;
20'b00000010000000001101:ColourData=12'h841;
20'b00000010010000001101:ColourData=12'h730;
20'b00000010100000001101:ColourData=12'h730;
20'b00000010110000001101:ColourData=12'h730;
20'b00000011000000001101:ColourData=12'h730;
20'b00000011010000001101:ColourData=12'h730;
20'b00000011100000001101:ColourData=12'h520;
20'b00000011110000001101:ColourData=12'h242;
20'b00000100000000001101:ColourData=12'h0D1;
20'b00000100010000001101:ColourData=12'h111;
20'b00000100100000001101:ColourData=12'h111;
20'b00000100110000001101:ColourData=12'h111;
20'b00000101000000001101:ColourData=12'h111;
20'b00000101010000001101:ColourData=12'h433;
20'b00000101100000001101:ColourData=12'hCA9;
20'b00000101110000001101:ColourData=12'hFCB;
20'b00000110000000001101:ColourData=12'hFCB;
20'b00000110010000001101:ColourData=12'hECA;
20'b00000110100000001101:ColourData=12'h876;
20'b00000110110000001101:ColourData=12'h101;
20'b00000111000000001101:ColourData=12'h060;
20'b00000111010000001101:ColourData=12'h0F0;
20'b00000111100000001101:ColourData=12'h0F0;
20'b00000111110000001101:ColourData=12'h6F6;
20'b00000000000000001110:ColourData=12'hD88;
20'b00000000010000001110:ColourData=12'h731;
20'b00000000100000001110:ColourData=12'h620;
20'b00000000110000001110:ColourData=12'h620;
20'b00000001000000001110:ColourData=12'h630;
20'b00000001010000001110:ColourData=12'h630;
20'b00000001100000001110:ColourData=12'h100;
20'b00000001110000001110:ColourData=12'hA55;
20'b00000010000000001110:ColourData=12'h731;
20'b00000010010000001110:ColourData=12'h620;
20'b00000010100000001110:ColourData=12'h630;
20'b00000010110000001110:ColourData=12'h630;
20'b00000011000000001110:ColourData=12'h630;
20'b00000011010000001110:ColourData=12'h520;
20'b00000011100000001110:ColourData=12'h000;
20'b00000011110000001110:ColourData=12'h242;
20'b00000100000000001110:ColourData=12'h0D1;
20'b00000100010000001110:ColourData=12'h140;
20'b00000100100000001110:ColourData=12'h111;
20'b00000100110000001110:ColourData=12'h111;
20'b00000101000000001110:ColourData=12'h111;
20'b00000101010000001110:ColourData=12'h101;
20'b00000101100000001110:ColourData=12'h343;
20'b00000101110000001110:ColourData=12'hAD8;
20'b00000110000000001110:ColourData=12'hBC8;
20'b00000110010000001110:ColourData=12'h876;
20'b00000110100000001110:ColourData=12'h101;
20'b00000110110000001110:ColourData=12'h111;
20'b00000111000000001110:ColourData=12'h080;
20'b00000111010000001110:ColourData=12'h0F0;
20'b00000111100000001110:ColourData=12'h0F0;
20'b00000111110000001110:ColourData=12'h6F6;
20'b00000000000000001111:ColourData=12'hA75;
20'b00000000010000001111:ColourData=12'h321;
20'b00000000100000001111:ColourData=12'h111;
20'b00000000110000001111:ColourData=12'h111;
20'b00000001000000001111:ColourData=12'h111;
20'b00000001010000001111:ColourData=12'h111;
20'b00000001100000001111:ColourData=12'h642;
20'b00000001110000001111:ColourData=12'hC77;
20'b00000010000000001111:ColourData=12'h322;
20'b00000010010000001111:ColourData=12'h111;
20'b00000010100000001111:ColourData=12'h111;
20'b00000010110000001111:ColourData=12'h111;
20'b00000011000000001111:ColourData=12'h111;
20'b00000011010000001111:ColourData=12'h111;
20'b00000011100000001111:ColourData=12'h111;
20'b00000011110000001111:ColourData=12'h774;
20'b00000100000000001111:ColourData=12'h0F0;
20'b00000100010000001111:ColourData=12'h0D0;
20'b00000100100000001111:ColourData=12'h141;
20'b00000100110000001111:ColourData=12'h141;
20'b00000101000000001111:ColourData=12'h041;
20'b00000101010000001111:ColourData=12'h131;
20'b00000101100000001111:ColourData=12'h350;
20'b00000101110000001111:ColourData=12'h2D0;
20'b00000110000000001111:ColourData=12'h390;
20'b00000110010000001111:ColourData=12'h331;
20'b00000110100000001111:ColourData=12'h041;
20'b00000110110000001111:ColourData=12'h080;
20'b00000111000000001111:ColourData=12'h0F0;
20'b00000111010000001111:ColourData=12'h0F0;
20'b00000111100000001111:ColourData=12'h0F0;
20'b00000111110000001111:ColourData=12'h6F6;
20'b00000000000000010000:ColourData=12'hEDD;
20'b00000000010000010000:ColourData=12'hDCC;
20'b00000000100000010000:ColourData=12'hDCC;
20'b00000000110000010000:ColourData=12'hDCC;
20'b00000001000000010000:ColourData=12'hDCC;
20'b00000001010000010000:ColourData=12'hDCC;
20'b00000001100000010000:ColourData=12'hDCC;
20'b00000001110000010000:ColourData=12'hDDD;
20'b00000010000000010000:ColourData=12'hDCC;
20'b00000010010000010000:ColourData=12'hDCC;
20'b00000010100000010000:ColourData=12'hDCC;
20'b00000010110000010000:ColourData=12'hDCC;
20'b00000011000000010000:ColourData=12'hDCC;
20'b00000011010000010000:ColourData=12'hDCC;
20'b00000011100000010000:ColourData=12'hDCC;
20'b00000011110000010000:ColourData=12'hBDB;
20'b00000100000000010000:ColourData=12'h0F0;
20'b00000100010000010000:ColourData=12'h0F0;
20'b00000100100000010000:ColourData=12'h0F0;
20'b00000100110000010000:ColourData=12'h0F0;
20'b00000101000000010000:ColourData=12'h0F0;
20'b00000101010000010000:ColourData=12'h5A0;
20'b00000101100000010000:ColourData=12'hD50;
20'b00000101110000010000:ColourData=12'hD50;
20'b00000110000000010000:ColourData=12'hD40;
20'b00000110010000010000:ColourData=12'hA70;
20'b00000110100000010000:ColourData=12'h1D0;
20'b00000110110000010000:ColourData=12'h0F0;
20'b00000111000000010000:ColourData=12'h0F0;
20'b00000111010000010000:ColourData=12'h0F0;
20'b00000111100000010000:ColourData=12'h0F0;
20'b00000111110000010000:ColourData=12'h6F6;
20'b00000000000000010001:ColourData=12'h944;
20'b00000000010000010001:ColourData=12'h811;
20'b00000000100000010001:ColourData=12'h812;
20'b00000000110000010001:ColourData=12'h812;
20'b00000001000000010001:ColourData=12'h812;
20'b00000001010000010001:ColourData=12'h812;
20'b00000001100000010001:ColourData=12'h711;
20'b00000001110000010001:ColourData=12'h211;
20'b00000010000000010001:ColourData=12'h711;
20'b00000010010000010001:ColourData=12'h812;
20'b00000010100000010001:ColourData=12'h812;
20'b00000010110000010001:ColourData=12'h812;
20'b00000011000000010001:ColourData=12'h812;
20'b00000011010000010001:ColourData=12'h812;
20'b00000011100000010001:ColourData=12'h711;
20'b00000011110000010001:ColourData=12'h353;
20'b00000100000000010001:ColourData=12'h0F0;
20'b00000100010000010001:ColourData=12'h0F0;
20'b00000100100000010001:ColourData=12'h0F0;
20'b00000100110000010001:ColourData=12'h0F0;
20'b00000101000000010001:ColourData=12'h5B0;
20'b00000101010000010001:ColourData=12'hD50;
20'b00000101100000010001:ColourData=12'hD40;
20'b00000101110000010001:ColourData=12'hD40;
20'b00000110000000010001:ColourData=12'hD40;
20'b00000110010000010001:ColourData=12'hE40;
20'b00000110100000010001:ColourData=12'hA70;
20'b00000110110000010001:ColourData=12'h1E0;
20'b00000111000000010001:ColourData=12'h0F0;
20'b00000111010000010001:ColourData=12'h0F0;
20'b00000111100000010001:ColourData=12'h0F0;
20'b00000111110000010001:ColourData=12'h6F6;
20'b00000000000000010010:ColourData=12'h823;
20'b00000000010000010010:ColourData=12'h500;
20'b00000000100000010010:ColourData=12'h600;
20'b00000000110000010010:ColourData=12'h600;
20'b00000001000000010010:ColourData=12'h600;
20'b00000001010000010010:ColourData=12'h600;
20'b00000001100000010010:ColourData=12'h500;
20'b00000001110000010010:ColourData=12'h000;
20'b00000010000000010010:ColourData=12'h500;
20'b00000010010000010010:ColourData=12'h600;
20'b00000010100000010010:ColourData=12'h600;
20'b00000010110000010010:ColourData=12'h600;
20'b00000011000000010010:ColourData=12'h600;
20'b00000011010000010010:ColourData=12'h600;
20'b00000011100000010010:ColourData=12'h500;
20'b00000011110000010010:ColourData=12'h232;
20'b00000100000000010010:ColourData=12'h0F0;
20'b00000100010000010010:ColourData=12'h0F0;
20'b00000100100000010010:ColourData=12'h0F0;
20'b00000100110000010010:ColourData=12'h5B0;
20'b00000101000000010010:ColourData=12'hD50;
20'b00000101010000010010:ColourData=12'hD40;
20'b00000101100000010010:ColourData=12'hD50;
20'b00000101110000010010:ColourData=12'hD50;
20'b00000110000000010010:ColourData=12'hD50;
20'b00000110010000010010:ColourData=12'hD50;
20'b00000110100000010010:ColourData=12'hE40;
20'b00000110110000010010:ColourData=12'hA70;
20'b00000111000000010010:ColourData=12'h1E0;
20'b00000111010000010010:ColourData=12'h0F0;
20'b00000111100000010010:ColourData=12'h0F0;
20'b00000111110000010010:ColourData=12'h6F6;
20'b00000000000000010011:ColourData=12'h433;
20'b00000000010000010011:ColourData=12'h000;
20'b00000000100000010011:ColourData=12'h000;
20'b00000000110000010011:ColourData=12'h000;
20'b00000001000000010011:ColourData=12'h000;
20'b00000001010000010011:ColourData=12'h000;
20'b00000001100000010011:ColourData=12'h000;
20'b00000001110000010011:ColourData=12'h000;
20'b00000010000000010011:ColourData=12'h000;
20'b00000010010000010011:ColourData=12'h000;
20'b00000010100000010011:ColourData=12'h000;
20'b00000010110000010011:ColourData=12'h000;
20'b00000011000000010011:ColourData=12'h000;
20'b00000011010000010011:ColourData=12'h000;
20'b00000011100000010011:ColourData=12'h000;
20'b00000011110000010011:ColourData=12'h242;
20'b00000100000000010011:ColourData=12'h0F0;
20'b00000100010000010011:ColourData=12'h0F0;
20'b00000100100000010011:ColourData=12'h4B0;
20'b00000100110000010011:ColourData=12'hA40;
20'b00000101000000010011:ColourData=12'hB40;
20'b00000101010000010011:ColourData=12'hE50;
20'b00000101100000010011:ColourData=12'hD50;
20'b00000101110000010011:ColourData=12'hD50;
20'b00000110000000010011:ColourData=12'hD50;
20'b00000110010000010011:ColourData=12'hE50;
20'b00000110100000010011:ColourData=12'hC40;
20'b00000110110000010011:ColourData=12'hA30;
20'b00000111000000010011:ColourData=12'h770;
20'b00000111010000010011:ColourData=12'h1E0;
20'b00000111100000010011:ColourData=12'h0F0;
20'b00000111110000010011:ColourData=12'h6F6;
20'b00000000000000010100:ColourData=12'h833;
20'b00000000010000010100:ColourData=12'h600;
20'b00000000100000010100:ColourData=12'h600;
20'b00000000110000010100:ColourData=12'h000;
20'b00000001000000010100:ColourData=12'h400;
20'b00000001010000010100:ColourData=12'h600;
20'b00000001100000010100:ColourData=12'h600;
20'b00000001110000010100:ColourData=12'h600;
20'b00000010000000010100:ColourData=12'h600;
20'b00000010010000010100:ColourData=12'h600;
20'b00000010100000010100:ColourData=12'h500;
20'b00000010110000010100:ColourData=12'h000;
20'b00000011000000010100:ColourData=12'h500;
20'b00000011010000010100:ColourData=12'h600;
20'b00000011100000010100:ColourData=12'h600;
20'b00000011110000010100:ColourData=12'h642;
20'b00000100000000010100:ColourData=12'h0F0;
20'b00000100010000010100:ColourData=12'h5B0;
20'b00000100100000010100:ColourData=12'hB40;
20'b00000100110000010100:ColourData=12'h421;
20'b00000101000000010100:ColourData=12'h642;
20'b00000101010000010100:ColourData=12'hB40;
20'b00000101100000010100:ColourData=12'hE50;
20'b00000101110000010100:ColourData=12'hE50;
20'b00000110000000010100:ColourData=12'hE50;
20'b00000110010000010100:ColourData=12'hD40;
20'b00000110100000010100:ColourData=12'h841;
20'b00000110110000010100:ColourData=12'h432;
20'b00000111000000010100:ColourData=12'h820;
20'b00000111010000010100:ColourData=12'h980;
20'b00000111100000010100:ColourData=12'h1E0;
20'b00000111110000010100:ColourData=12'h6F6;
20'b00000000000000010101:ColourData=12'h933;
20'b00000000010000010101:ColourData=12'h700;
20'b00000000100000010101:ColourData=12'h700;
20'b00000000110000010101:ColourData=12'h100;
20'b00000001000000010101:ColourData=12'h500;
20'b00000001010000010101:ColourData=12'h700;
20'b00000001100000010101:ColourData=12'h700;
20'b00000001110000010101:ColourData=12'h700;
20'b00000010000000010101:ColourData=12'h700;
20'b00000010010000010101:ColourData=12'h700;
20'b00000010100000010101:ColourData=12'h600;
20'b00000010110000010101:ColourData=12'h100;
20'b00000011000000010101:ColourData=12'h600;
20'b00000011010000010101:ColourData=12'h700;
20'b00000011100000010101:ColourData=12'h700;
20'b00000011110000010101:ColourData=12'h742;
20'b00000100000000010101:ColourData=12'h2D0;
20'b00000100010000010101:ColourData=12'hD50;
20'b00000100100000010101:ColourData=12'hD40;
20'b00000100110000010101:ColourData=12'hE73;
20'b00000101000000010101:ColourData=12'hB98;
20'b00000101010000010101:ColourData=12'h321;
20'b00000101100000010101:ColourData=12'hA30;
20'b00000101110000010101:ColourData=12'hA40;
20'b00000110000000010101:ColourData=12'hA40;
20'b00000110010000010101:ColourData=12'h720;
20'b00000110100000010101:ColourData=12'h554;
20'b00000110110000010101:ColourData=12'hEA7;
20'b00000111000000010101:ColourData=12'hD40;
20'b00000111010000010101:ColourData=12'hE40;
20'b00000111100000010101:ColourData=12'h790;
20'b00000111110000010101:ColourData=12'h5F6;
20'b00000000000000010110:ColourData=12'h833;
20'b00000000010000010110:ColourData=12'h600;
20'b00000000100000010110:ColourData=12'h600;
20'b00000000110000010110:ColourData=12'h000;
20'b00000001000000010110:ColourData=12'h400;
20'b00000001010000010110:ColourData=12'h600;
20'b00000001100000010110:ColourData=12'h600;
20'b00000001110000010110:ColourData=12'h600;
20'b00000010000000010110:ColourData=12'h600;
20'b00000010010000010110:ColourData=12'h600;
20'b00000010100000010110:ColourData=12'h500;
20'b00000010110000010110:ColourData=12'h000;
20'b00000011000000010110:ColourData=12'h500;
20'b00000011010000010110:ColourData=12'h600;
20'b00000011100000010110:ColourData=12'h600;
20'b00000011110000010110:ColourData=12'h742;
20'b00000100000000010110:ColourData=12'h5B1;
20'b00000100010000010110:ColourData=12'hD50;
20'b00000100100000010110:ColourData=12'hD40;
20'b00000100110000010110:ColourData=12'hE73;
20'b00000101000000010110:ColourData=12'hB98;
20'b00000101010000010110:ColourData=12'h222;
20'b00000101100000010110:ColourData=12'h432;
20'b00000101110000010110:ColourData=12'h421;
20'b00000110000000010110:ColourData=12'h422;
20'b00000110010000010110:ColourData=12'h322;
20'b00000110100000010110:ColourData=12'h554;
20'b00000110110000010110:ColourData=12'hEA7;
20'b00000111000000010110:ColourData=12'hD40;
20'b00000111010000010110:ColourData=12'hE40;
20'b00000111100000010110:ColourData=12'h970;
20'b00000111110000010110:ColourData=12'h7E6;
20'b00000000000000010111:ColourData=12'h433;
20'b00000000010000010111:ColourData=12'h000;
20'b00000000100000010111:ColourData=12'h000;
20'b00000000110000010111:ColourData=12'h000;
20'b00000001000000010111:ColourData=12'h000;
20'b00000001010000010111:ColourData=12'h000;
20'b00000001100000010111:ColourData=12'h000;
20'b00000001110000010111:ColourData=12'h000;
20'b00000010000000010111:ColourData=12'h000;
20'b00000010010000010111:ColourData=12'h000;
20'b00000010100000010111:ColourData=12'h000;
20'b00000010110000010111:ColourData=12'h000;
20'b00000011000000010111:ColourData=12'h000;
20'b00000011010000010111:ColourData=12'h000;
20'b00000011100000010111:ColourData=12'h000;
20'b00000011110000010111:ColourData=12'h422;
20'b00000100000000010111:ColourData=12'hD51;
20'b00000100010000010111:ColourData=12'hD40;
20'b00000100100000010111:ColourData=12'hD40;
20'b00000100110000010111:ColourData=12'hE73;
20'b00000101000000010111:ColourData=12'hCA9;
20'b00000101010000010111:ColourData=12'h766;
20'b00000101100000010111:ColourData=12'hEA8;
20'b00000101110000010111:ColourData=12'hD40;
20'b00000110000000010111:ColourData=12'hE73;
20'b00000110010000010111:ColourData=12'hB98;
20'b00000110100000010111:ColourData=12'h776;
20'b00000110110000010111:ColourData=12'hEA7;
20'b00000111000000010111:ColourData=12'hD40;
20'b00000111010000010111:ColourData=12'hD50;
20'b00000111100000010111:ColourData=12'hD40;
20'b00000111110000010111:ColourData=12'hE96;
20'b00000000000000011000:ColourData=12'h833;
20'b00000000010000011000:ColourData=12'h600;
20'b00000000100000011000:ColourData=12'h600;
20'b00000000110000011000:ColourData=12'h600;
20'b00000001000000011000:ColourData=12'h600;
20'b00000001010000011000:ColourData=12'h600;
20'b00000001100000011000:ColourData=12'h500;
20'b00000001110000011000:ColourData=12'h000;
20'b00000010000000011000:ColourData=12'h500;
20'b00000010010000011000:ColourData=12'h600;
20'b00000010100000011000:ColourData=12'h600;
20'b00000010110000011000:ColourData=12'h600;
20'b00000011000000011000:ColourData=12'h600;
20'b00000011010000011000:ColourData=12'h600;
20'b00000011100000011000:ColourData=12'h500;
20'b00000011110000011000:ColourData=12'h422;
20'b00000100000000011000:ColourData=12'hE51;
20'b00000100010000011000:ColourData=12'hD40;
20'b00000100100000011000:ColourData=12'hD40;
20'b00000100110000011000:ColourData=12'hD62;
20'b00000101000000011000:ColourData=12'hEA8;
20'b00000101010000011000:ColourData=12'hEA8;
20'b00000101100000011000:ColourData=12'hE96;
20'b00000101110000011000:ColourData=12'hD40;
20'b00000110000000011000:ColourData=12'hE62;
20'b00000110010000011000:ColourData=12'hEA8;
20'b00000110100000011000:ColourData=12'hEB8;
20'b00000110110000011000:ColourData=12'hE85;
20'b00000111000000011000:ColourData=12'hD40;
20'b00000111010000011000:ColourData=12'hD50;
20'b00000111100000011000:ColourData=12'hD40;
20'b00000111110000011000:ColourData=12'hE96;
20'b00000000000000011001:ColourData=12'h933;
20'b00000000010000011001:ColourData=12'h700;
20'b00000000100000011001:ColourData=12'h700;
20'b00000000110000011001:ColourData=12'h700;
20'b00000001000000011001:ColourData=12'h700;
20'b00000001010000011001:ColourData=12'h700;
20'b00000001100000011001:ColourData=12'h600;
20'b00000001110000011001:ColourData=12'h100;
20'b00000010000000011001:ColourData=12'h600;
20'b00000010010000011001:ColourData=12'h700;
20'b00000010100000011001:ColourData=12'h700;
20'b00000010110000011001:ColourData=12'h700;
20'b00000011000000011001:ColourData=12'h700;
20'b00000011010000011001:ColourData=12'h700;
20'b00000011100000011001:ColourData=12'h600;
20'b00000011110000011001:ColourData=12'h332;
20'b00000100000000011001:ColourData=12'hB71;
20'b00000100010000011001:ColourData=12'hE40;
20'b00000100100000011001:ColourData=12'hE40;
20'b00000100110000011001:ColourData=12'hE40;
20'b00000101000000011001:ColourData=12'hD51;
20'b00000101010000011001:ColourData=12'hE63;
20'b00000101100000011001:ColourData=12'hE62;
20'b00000101110000011001:ColourData=12'hE62;
20'b00000110000000011001:ColourData=12'hD62;
20'b00000110010000011001:ColourData=12'hE63;
20'b00000110100000011001:ColourData=12'hD62;
20'b00000110110000011001:ColourData=12'hD40;
20'b00000111000000011001:ColourData=12'hE40;
20'b00000111010000011001:ColourData=12'hE40;
20'b00000111100000011001:ColourData=12'hC50;
20'b00000111110000011001:ColourData=12'hCA6;
20'b00000000000000011010:ColourData=12'h833;
20'b00000000010000011010:ColourData=12'h600;
20'b00000000100000011010:ColourData=12'h600;
20'b00000000110000011010:ColourData=12'h600;
20'b00000001000000011010:ColourData=12'h600;
20'b00000001010000011010:ColourData=12'h600;
20'b00000001100000011010:ColourData=12'h500;
20'b00000001110000011010:ColourData=12'h000;
20'b00000010000000011010:ColourData=12'h500;
20'b00000010010000011010:ColourData=12'h600;
20'b00000010100000011010:ColourData=12'h600;
20'b00000010110000011010:ColourData=12'h600;
20'b00000011000000011010:ColourData=12'h600;
20'b00000011010000011010:ColourData=12'h600;
20'b00000011100000011010:ColourData=12'h500;
20'b00000011110000011010:ColourData=12'h242;
20'b00000100000000011010:ColourData=12'h2E0;
20'b00000100010000011010:ColourData=12'hA70;
20'b00000100100000011010:ColourData=12'hA70;
20'b00000100110000011010:ColourData=12'hB70;
20'b00000101000000011010:ColourData=12'hE84;
20'b00000101010000011010:ColourData=12'hECA;
20'b00000101100000011010:ColourData=12'hECA;
20'b00000101110000011010:ColourData=12'hECA;
20'b00000110000000011010:ColourData=12'hECA;
20'b00000110010000011010:ColourData=12'hECA;
20'b00000110100000011010:ColourData=12'hEA8;
20'b00000110110000011010:ColourData=12'hC71;
20'b00000111000000011010:ColourData=12'hA70;
20'b00000111010000011010:ColourData=12'hA70;
20'b00000111100000011010:ColourData=12'h5A0;
20'b00000111110000011010:ColourData=12'h6F6;
20'b00000000000000011011:ColourData=12'h433;
20'b00000000010000011011:ColourData=12'h000;
20'b00000000100000011011:ColourData=12'h000;
20'b00000000110000011011:ColourData=12'h000;
20'b00000001000000011011:ColourData=12'h000;
20'b00000001010000011011:ColourData=12'h000;
20'b00000001100000011011:ColourData=12'h000;
20'b00000001110000011011:ColourData=12'h000;
20'b00000010000000011011:ColourData=12'h000;
20'b00000010010000011011:ColourData=12'h000;
20'b00000010100000011011:ColourData=12'h000;
20'b00000010110000011011:ColourData=12'h000;
20'b00000011000000011011:ColourData=12'h000;
20'b00000011010000011011:ColourData=12'h000;
20'b00000011100000011011:ColourData=12'h000;
20'b00000011110000011011:ColourData=12'h242;
20'b00000100000000011011:ColourData=12'h0F0;
20'b00000100010000011011:ColourData=12'h0F0;
20'b00000100100000011011:ColourData=12'h0F0;
20'b00000100110000011011:ColourData=12'h3F2;
20'b00000101000000011011:ColourData=12'hECA;
20'b00000101010000011011:ColourData=12'hECA;
20'b00000101100000011011:ColourData=12'hECA;
20'b00000101110000011011:ColourData=12'hECA;
20'b00000110000000011011:ColourData=12'hECA;
20'b00000110010000011011:ColourData=12'hECA;
20'b00000110100000011011:ColourData=12'hFDB;
20'b00000110110000011011:ColourData=12'hAC7;
20'b00000111000000011011:ColourData=12'h0B0;
20'b00000111010000011011:ColourData=12'h0D0;
20'b00000111100000011011:ColourData=12'h0F0;
20'b00000111110000011011:ColourData=12'h6F6;
20'b00000000000000011100:ColourData=12'h833;
20'b00000000010000011100:ColourData=12'h600;
20'b00000000100000011100:ColourData=12'h600;
20'b00000000110000011100:ColourData=12'h000;
20'b00000001000000011100:ColourData=12'h400;
20'b00000001010000011100:ColourData=12'h600;
20'b00000001100000011100:ColourData=12'h600;
20'b00000001110000011100:ColourData=12'h600;
20'b00000010000000011100:ColourData=12'h600;
20'b00000010010000011100:ColourData=12'h600;
20'b00000010100000011100:ColourData=12'h500;
20'b00000010110000011100:ColourData=12'h000;
20'b00000011000000011100:ColourData=12'h500;
20'b00000011010000011100:ColourData=12'h600;
20'b00000011100000011100:ColourData=12'h600;
20'b00000011110000011100:ColourData=12'h742;
20'b00000100000000011100:ColourData=12'h0F0;
20'b00000100010000011100:ColourData=12'h0F0;
20'b00000100100000011100:ColourData=12'h0E0;
20'b00000100110000011100:ColourData=12'h2B1;
20'b00000101000000011100:ColourData=12'hCA9;
20'b00000101010000011100:ColourData=12'hFCA;
20'b00000101100000011100:ColourData=12'hECA;
20'b00000101110000011100:ColourData=12'hECA;
20'b00000110000000011100:ColourData=12'hECA;
20'b00000110010000011100:ColourData=12'hECA;
20'b00000110100000011100:ColourData=12'hCA8;
20'b00000110110000011100:ColourData=12'h876;
20'b00000111000000011100:ColourData=12'h111;
20'b00000111010000011100:ColourData=12'h050;
20'b00000111100000011100:ColourData=12'h0D0;
20'b00000111110000011100:ColourData=12'h6F6;
20'b00000000000000011101:ColourData=12'h933;
20'b00000000010000011101:ColourData=12'h700;
20'b00000000100000011101:ColourData=12'h700;
20'b00000000110000011101:ColourData=12'h100;
20'b00000001000000011101:ColourData=12'h500;
20'b00000001010000011101:ColourData=12'h700;
20'b00000001100000011101:ColourData=12'h700;
20'b00000001110000011101:ColourData=12'h700;
20'b00000010000000011101:ColourData=12'h700;
20'b00000010010000011101:ColourData=12'h700;
20'b00000010100000011101:ColourData=12'h600;
20'b00000010110000011101:ColourData=12'h100;
20'b00000011000000011101:ColourData=12'h600;
20'b00000011010000011101:ColourData=12'h700;
20'b00000011100000011101:ColourData=12'h700;
20'b00000011110000011101:ColourData=12'h742;
20'b00000100000000011101:ColourData=12'h0F0;
20'b00000100010000011101:ColourData=12'h0F0;
20'b00000100100000011101:ColourData=12'h0C0;
20'b00000100110000011101:ColourData=12'h111;
20'b00000101000000011101:ColourData=12'h433;
20'b00000101010000011101:ColourData=12'hCA9;
20'b00000101100000011101:ColourData=12'hFDB;
20'b00000101110000011101:ColourData=12'hFCB;
20'b00000110000000011101:ColourData=12'hECA;
20'b00000110010000011101:ColourData=12'h876;
20'b00000110100000011101:ColourData=12'h111;
20'b00000110110000011101:ColourData=12'h111;
20'b00000111000000011101:ColourData=12'h111;
20'b00000111010000011101:ColourData=12'h101;
20'b00000111100000011101:ColourData=12'h060;
20'b00000111110000011101:ColourData=12'h6F6;
20'b00000000000000011110:ColourData=12'h823;
20'b00000000010000011110:ColourData=12'h600;
20'b00000000100000011110:ColourData=12'h600;
20'b00000000110000011110:ColourData=12'h000;
20'b00000001000000011110:ColourData=12'h400;
20'b00000001010000011110:ColourData=12'h600;
20'b00000001100000011110:ColourData=12'h600;
20'b00000001110000011110:ColourData=12'h600;
20'b00000010000000011110:ColourData=12'h600;
20'b00000010010000011110:ColourData=12'h600;
20'b00000010100000011110:ColourData=12'h500;
20'b00000010110000011110:ColourData=12'h000;
20'b00000011000000011110:ColourData=12'h500;
20'b00000011010000011110:ColourData=12'h600;
20'b00000011100000011110:ColourData=12'h600;
20'b00000011110000011110:ColourData=12'h742;
20'b00000100000000011110:ColourData=12'h0F0;
20'b00000100010000011110:ColourData=12'h0F0;
20'b00000100100000011110:ColourData=12'h0D0;
20'b00000100110000011110:ColourData=12'h131;
20'b00000101000000011110:ColourData=12'h101;
20'b00000101010000011110:ColourData=12'h433;
20'b00000101100000011110:ColourData=12'hBA8;
20'b00000101110000011110:ColourData=12'hBD8;
20'b00000110000000011110:ColourData=12'h896;
20'b00000110010000011110:ColourData=12'h111;
20'b00000110100000011110:ColourData=12'h111;
20'b00000110110000011110:ColourData=12'h111;
20'b00000111000000011110:ColourData=12'h111;
20'b00000111010000011110:ColourData=12'h121;
20'b00000111100000011110:ColourData=12'h080;
20'b00000111110000011110:ColourData=12'h6F6;
20'b00000000000000011111:ColourData=12'h433;
20'b00000000010000011111:ColourData=12'h100;
20'b00000000100000011111:ColourData=12'h100;
20'b00000000110000011111:ColourData=12'h000;
20'b00000001000000011111:ColourData=12'h100;
20'b00000001010000011111:ColourData=12'h100;
20'b00000001100000011111:ColourData=12'h100;
20'b00000001110000011111:ColourData=12'h100;
20'b00000010000000011111:ColourData=12'h100;
20'b00000010010000011111:ColourData=12'h100;
20'b00000010100000011111:ColourData=12'h100;
20'b00000010110000011111:ColourData=12'h000;
20'b00000011000000011111:ColourData=12'h100;
20'b00000011010000011111:ColourData=12'h100;
20'b00000011100000011111:ColourData=12'h100;
20'b00000011110000011111:ColourData=12'h242;
20'b00000100000000011111:ColourData=12'h0F0;
20'b00000100010000011111:ColourData=12'h0F0;
20'b00000100100000011111:ColourData=12'h0F0;
20'b00000100110000011111:ColourData=12'h0C0;
20'b00000101000000011111:ColourData=12'h141;
20'b00000101010000011111:ColourData=12'h141;
20'b00000101100000011111:ColourData=12'h070;
20'b00000101110000011111:ColourData=12'h0F0;
20'b00000110000000011111:ColourData=12'h0C0;
20'b00000110010000011111:ColourData=12'h141;
20'b00000110100000011111:ColourData=12'h141;
20'b00000110110000011111:ColourData=12'h141;
20'b00000111000000011111:ColourData=12'h141;
20'b00000111010000011111:ColourData=12'h080;
20'b00000111100000011111:ColourData=12'h0F0;
20'b00000111110000011111:ColourData=12'h6F6;
20'b00000000000000100000:ColourData=12'h864;
20'b00000000010000100000:ColourData=12'h954;
20'b00000000100000100000:ColourData=12'hB66;
20'b00000000110000100000:ColourData=12'hB66;
20'b00000001000000100000:ColourData=12'hB66;
20'b00000001010000100000:ColourData=12'hB66;
20'b00000001100000100000:ColourData=12'hB66;
20'b00000001110000100000:ColourData=12'hB66;
20'b00000010000000100000:ColourData=12'hB66;
20'b00000010010000100000:ColourData=12'hB66;
20'b00000010100000100000:ColourData=12'hB66;
20'b00000010110000100000:ColourData=12'hB66;
20'b00000011000000100000:ColourData=12'hB66;
20'b00000011010000100000:ColourData=12'hB66;
20'b00000011100000100000:ColourData=12'h845;
20'b00000011110000100000:ColourData=12'h342;
20'b00000100000000100000:ColourData=12'h0F0;
20'b00000100010000100000:ColourData=12'h0F0;
20'b00000100100000100000:ColourData=12'h0F0;
20'b00000100110000100000:ColourData=12'h0F0;
20'b00000101000000100000:ColourData=12'h0F0;
20'b00000101010000100000:ColourData=12'h0F0;
20'b00000101100000100000:ColourData=12'h0F0;
20'b00000101110000100000:ColourData=12'h0F0;
20'b00000110000000100000:ColourData=12'h0F0;
20'b00000110010000100000:ColourData=12'h0F0;
20'b00000110100000100000:ColourData=12'h0F0;
20'b00000110110000100000:ColourData=12'h0F0;
20'b00000111000000100000:ColourData=12'h0F0;
20'b00000111010000100000:ColourData=12'h0F0;
20'b00000111100000100000:ColourData=12'h0F0;
20'b00000111110000100000:ColourData=12'h6F6;
20'b00000000000000100001:ColourData=12'hD88;
20'b00000000010000100001:ColourData=12'h942;
20'b00000000100000100001:ColourData=12'hB65;
20'b00000000110000100001:ColourData=12'hD77;
20'b00000001000000100001:ColourData=12'hD77;
20'b00000001010000100001:ColourData=12'hD77;
20'b00000001100000100001:ColourData=12'hD77;
20'b00000001110000100001:ColourData=12'hD77;
20'b00000010000000100001:ColourData=12'hD77;
20'b00000010010000100001:ColourData=12'hD77;
20'b00000010100000100001:ColourData=12'hD77;
20'b00000010110000100001:ColourData=12'hD77;
20'b00000011000000100001:ColourData=12'hD77;
20'b00000011010000100001:ColourData=12'hA66;
20'b00000011100000100001:ColourData=12'h100;
20'b00000011110000100001:ColourData=12'h242;
20'b00000100000000100001:ColourData=12'h0F0;
20'b00000100010000100001:ColourData=12'h0F0;
20'b00000100100000100001:ColourData=12'h0F0;
20'b00000100110000100001:ColourData=12'h0F0;
20'b00000101000000100001:ColourData=12'h0F0;
20'b00000101010000100001:ColourData=12'h0F0;
20'b00000101100000100001:ColourData=12'h0F0;
20'b00000101110000100001:ColourData=12'h0F0;
20'b00000110000000100001:ColourData=12'h0F0;
20'b00000110010000100001:ColourData=12'h0F0;
20'b00000110100000100001:ColourData=12'h0F0;
20'b00000110110000100001:ColourData=12'h0F0;
20'b00000111000000100001:ColourData=12'h0F0;
20'b00000111010000100001:ColourData=12'h0F0;
20'b00000111100000100001:ColourData=12'h0F0;
20'b00000111110000100001:ColourData=12'h6F6;
20'b00000000000000100010:ColourData=12'hD99;
20'b00000000010000100010:ColourData=12'hC66;
20'b00000000100000100010:ColourData=12'h942;
20'b00000000110000100010:ColourData=12'hB65;
20'b00000001000000100010:ColourData=12'hD77;
20'b00000001010000100010:ColourData=12'hD77;
20'b00000001100000100010:ColourData=12'hD77;
20'b00000001110000100010:ColourData=12'hD77;
20'b00000010000000100010:ColourData=12'hD77;
20'b00000010010000100010:ColourData=12'hD77;
20'b00000010100000100010:ColourData=12'hD77;
20'b00000010110000100010:ColourData=12'hD77;
20'b00000011000000100010:ColourData=12'hA66;
20'b00000011010000100010:ColourData=12'h100;
20'b00000011100000100010:ColourData=12'h000;
20'b00000011110000100010:ColourData=12'h242;
20'b00000100000000100010:ColourData=12'h0F0;
20'b00000100010000100010:ColourData=12'h0F0;
20'b00000100100000100010:ColourData=12'h0F0;
20'b00000100110000100010:ColourData=12'h0F0;
20'b00000101000000100010:ColourData=12'h0F0;
20'b00000101010000100010:ColourData=12'h0F0;
20'b00000101100000100010:ColourData=12'h0F0;
20'b00000101110000100010:ColourData=12'h0F0;
20'b00000110000000100010:ColourData=12'h0F0;
20'b00000110010000100010:ColourData=12'h0F0;
20'b00000110100000100010:ColourData=12'h0F0;
20'b00000110110000100010:ColourData=12'h0F0;
20'b00000111000000100010:ColourData=12'h0F0;
20'b00000111010000100010:ColourData=12'h0F0;
20'b00000111100000100010:ColourData=12'h0F0;
20'b00000111110000100010:ColourData=12'h6F6;
20'b00000000000000100011:ColourData=12'hD99;
20'b00000000010000100011:ColourData=12'hD77;
20'b00000000100000100011:ColourData=12'hC66;
20'b00000000110000100011:ColourData=12'h942;
20'b00000001000000100011:ColourData=12'hB65;
20'b00000001010000100011:ColourData=12'hC76;
20'b00000001100000100011:ColourData=12'hC66;
20'b00000001110000100011:ColourData=12'hC66;
20'b00000010000000100011:ColourData=12'hC66;
20'b00000010010000100011:ColourData=12'hC66;
20'b00000010100000100011:ColourData=12'hC76;
20'b00000010110000100011:ColourData=12'hB66;
20'b00000011000000100011:ColourData=12'h100;
20'b00000011010000100011:ColourData=12'h000;
20'b00000011100000100011:ColourData=12'h000;
20'b00000011110000100011:ColourData=12'h242;
20'b00000100000000100011:ColourData=12'h0F0;
20'b00000100010000100011:ColourData=12'h0F0;
20'b00000100100000100011:ColourData=12'h0F0;
20'b00000100110000100011:ColourData=12'h0F0;
20'b00000101000000100011:ColourData=12'h0F0;
20'b00000101010000100011:ColourData=12'h0F0;
20'b00000101100000100011:ColourData=12'h0F0;
20'b00000101110000100011:ColourData=12'h0F0;
20'b00000110000000100011:ColourData=12'h0F0;
20'b00000110010000100011:ColourData=12'h0F0;
20'b00000110100000100011:ColourData=12'h0F0;
20'b00000110110000100011:ColourData=12'h0F0;
20'b00000111000000100011:ColourData=12'h0F0;
20'b00000111010000100011:ColourData=12'h0F0;
20'b00000111100000100011:ColourData=12'h0F0;
20'b00000111110000100011:ColourData=12'h6F6;
20'b00000000000000100100:ColourData=12'hD99;
20'b00000000010000100100:ColourData=12'hD77;
20'b00000000100000100100:ColourData=12'hD77;
20'b00000000110000100100:ColourData=12'hC66;
20'b00000001000000100100:ColourData=12'h842;
20'b00000001010000100100:ColourData=12'h731;
20'b00000001100000100100:ColourData=12'h731;
20'b00000001110000100100:ColourData=12'h731;
20'b00000010000000100100:ColourData=12'h731;
20'b00000010010000100100:ColourData=12'h731;
20'b00000010100000100100:ColourData=12'h741;
20'b00000010110000100100:ColourData=12'h730;
20'b00000011000000100100:ColourData=12'h000;
20'b00000011010000100100:ColourData=12'h000;
20'b00000011100000100100:ColourData=12'h000;
20'b00000011110000100100:ColourData=12'h242;
20'b00000100000000100100:ColourData=12'h0F0;
20'b00000100010000100100:ColourData=12'h0F0;
20'b00000100100000100100:ColourData=12'h0F0;
20'b00000100110000100100:ColourData=12'h0F0;
20'b00000101000000100100:ColourData=12'h0F0;
20'b00000101010000100100:ColourData=12'h0F0;
20'b00000101100000100100:ColourData=12'h0F0;
20'b00000101110000100100:ColourData=12'h0F0;
20'b00000110000000100100:ColourData=12'h0F0;
20'b00000110010000100100:ColourData=12'h0F0;
20'b00000110100000100100:ColourData=12'h0F0;
20'b00000110110000100100:ColourData=12'h0F0;
20'b00000111000000100100:ColourData=12'h0F0;
20'b00000111010000100100:ColourData=12'h0F0;
20'b00000111100000100100:ColourData=12'h0F0;
20'b00000111110000100100:ColourData=12'h6F6;
20'b00000000000000100101:ColourData=12'hD99;
20'b00000000010000100101:ColourData=12'hD77;
20'b00000000100000100101:ColourData=12'hD77;
20'b00000000110000100101:ColourData=12'hC77;
20'b00000001000000100101:ColourData=12'h841;
20'b00000001010000100101:ColourData=12'h730;
20'b00000001100000100101:ColourData=12'h730;
20'b00000001110000100101:ColourData=12'h730;
20'b00000010000000100101:ColourData=12'h730;
20'b00000010010000100101:ColourData=12'h730;
20'b00000010100000100101:ColourData=12'h730;
20'b00000010110000100101:ColourData=12'h630;
20'b00000011000000100101:ColourData=12'h000;
20'b00000011010000100101:ColourData=12'h000;
20'b00000011100000100101:ColourData=12'h000;
20'b00000011110000100101:ColourData=12'h242;
20'b00000100000000100101:ColourData=12'h0F0;
20'b00000100010000100101:ColourData=12'h0F0;
20'b00000100100000100101:ColourData=12'h0F0;
20'b00000100110000100101:ColourData=12'h0F0;
20'b00000101000000100101:ColourData=12'h0F0;
20'b00000101010000100101:ColourData=12'h0F0;
20'b00000101100000100101:ColourData=12'h0F0;
20'b00000101110000100101:ColourData=12'h0F0;
20'b00000110000000100101:ColourData=12'h0F0;
20'b00000110010000100101:ColourData=12'h0F0;
20'b00000110100000100101:ColourData=12'h0F0;
20'b00000110110000100101:ColourData=12'h0F0;
20'b00000111000000100101:ColourData=12'h0F0;
20'b00000111010000100101:ColourData=12'h0F0;
20'b00000111100000100101:ColourData=12'h0F0;
20'b00000111110000100101:ColourData=12'h6F6;
20'b00000000000000100110:ColourData=12'hD99;
20'b00000000010000100110:ColourData=12'hD77;
20'b00000000100000100110:ColourData=12'hD77;
20'b00000000110000100110:ColourData=12'hC77;
20'b00000001000000100110:ColourData=12'h841;
20'b00000001010000100110:ColourData=12'h730;
20'b00000001100000100110:ColourData=12'h730;
20'b00000001110000100110:ColourData=12'h730;
20'b00000010000000100110:ColourData=12'h730;
20'b00000010010000100110:ColourData=12'h730;
20'b00000010100000100110:ColourData=12'h730;
20'b00000010110000100110:ColourData=12'h630;
20'b00000011000000100110:ColourData=12'h000;
20'b00000011010000100110:ColourData=12'h000;
20'b00000011100000100110:ColourData=12'h000;
20'b00000011110000100110:ColourData=12'h242;
20'b00000100000000100110:ColourData=12'h0F0;
20'b00000100010000100110:ColourData=12'h0F0;
20'b00000100100000100110:ColourData=12'h0F0;
20'b00000100110000100110:ColourData=12'h0F0;
20'b00000101000000100110:ColourData=12'h0F0;
20'b00000101010000100110:ColourData=12'h0F0;
20'b00000101100000100110:ColourData=12'h0F0;
20'b00000101110000100110:ColourData=12'h0F0;
20'b00000110000000100110:ColourData=12'h0F0;
20'b00000110010000100110:ColourData=12'h0F0;
20'b00000110100000100110:ColourData=12'h0F0;
20'b00000110110000100110:ColourData=12'h0F0;
20'b00000111000000100110:ColourData=12'h0F0;
20'b00000111010000100110:ColourData=12'h0F0;
20'b00000111100000100110:ColourData=12'h0F0;
20'b00000111110000100110:ColourData=12'h6F6;
20'b00000000000000100111:ColourData=12'hD99;
20'b00000000010000100111:ColourData=12'hD77;
20'b00000000100000100111:ColourData=12'hD77;
20'b00000000110000100111:ColourData=12'hC77;
20'b00000001000000100111:ColourData=12'h841;
20'b00000001010000100111:ColourData=12'h730;
20'b00000001100000100111:ColourData=12'h730;
20'b00000001110000100111:ColourData=12'h730;
20'b00000010000000100111:ColourData=12'h730;
20'b00000010010000100111:ColourData=12'h730;
20'b00000010100000100111:ColourData=12'h730;
20'b00000010110000100111:ColourData=12'h630;
20'b00000011000000100111:ColourData=12'h000;
20'b00000011010000100111:ColourData=12'h000;
20'b00000011100000100111:ColourData=12'h000;
20'b00000011110000100111:ColourData=12'h242;
20'b00000100000000100111:ColourData=12'h0F0;
20'b00000100010000100111:ColourData=12'h0F0;
20'b00000100100000100111:ColourData=12'h0F0;
20'b00000100110000100111:ColourData=12'h0F0;
20'b00000101000000100111:ColourData=12'h0F0;
20'b00000101010000100111:ColourData=12'h0F0;
20'b00000101100000100111:ColourData=12'h2D0;
20'b00000101110000100111:ColourData=12'h2D0;
20'b00000110000000100111:ColourData=12'h2C0;
20'b00000110010000100111:ColourData=12'h1D0;
20'b00000110100000100111:ColourData=12'h0F0;
20'b00000110110000100111:ColourData=12'h0F0;
20'b00000111000000100111:ColourData=12'h0F0;
20'b00000111010000100111:ColourData=12'h0F0;
20'b00000111100000100111:ColourData=12'h0F0;
20'b00000111110000100111:ColourData=12'h6F6;
20'b00000000000000101000:ColourData=12'hD99;
20'b00000000010000101000:ColourData=12'hD77;
20'b00000000100000101000:ColourData=12'hD77;
20'b00000000110000101000:ColourData=12'hC77;
20'b00000001000000101000:ColourData=12'h841;
20'b00000001010000101000:ColourData=12'h730;
20'b00000001100000101000:ColourData=12'h730;
20'b00000001110000101000:ColourData=12'h730;
20'b00000010000000101000:ColourData=12'h730;
20'b00000010010000101000:ColourData=12'h730;
20'b00000010100000101000:ColourData=12'h730;
20'b00000010110000101000:ColourData=12'h630;
20'b00000011000000101000:ColourData=12'h000;
20'b00000011010000101000:ColourData=12'h000;
20'b00000011100000101000:ColourData=12'h000;
20'b00000011110000101000:ColourData=12'h242;
20'b00000100000000101000:ColourData=12'h0F0;
20'b00000100010000101000:ColourData=12'h0F0;
20'b00000100100000101000:ColourData=12'h0F0;
20'b00000100110000101000:ColourData=12'h3D0;
20'b00000101000000101000:ColourData=12'h3D0;
20'b00000101010000101000:ColourData=12'h5B0;
20'b00000101100000101000:ColourData=12'hD50;
20'b00000101110000101000:ColourData=12'hD50;
20'b00000110000000101000:ColourData=12'hD40;
20'b00000110010000101000:ColourData=12'hA70;
20'b00000110100000101000:ColourData=12'h3D0;
20'b00000110110000101000:ColourData=12'h3D0;
20'b00000111000000101000:ColourData=12'h1E0;
20'b00000111010000101000:ColourData=12'h0F0;
20'b00000111100000101000:ColourData=12'h0F0;
20'b00000111110000101000:ColourData=12'h6F6;
20'b00000000000000101001:ColourData=12'hD99;
20'b00000000010000101001:ColourData=12'hD77;
20'b00000000100000101001:ColourData=12'hD77;
20'b00000000110000101001:ColourData=12'hC77;
20'b00000001000000101001:ColourData=12'h841;
20'b00000001010000101001:ColourData=12'h730;
20'b00000001100000101001:ColourData=12'h730;
20'b00000001110000101001:ColourData=12'h730;
20'b00000010000000101001:ColourData=12'h730;
20'b00000010010000101001:ColourData=12'h730;
20'b00000010100000101001:ColourData=12'h730;
20'b00000010110000101001:ColourData=12'h630;
20'b00000011000000101001:ColourData=12'h000;
20'b00000011010000101001:ColourData=12'h000;
20'b00000011100000101001:ColourData=12'h000;
20'b00000011110000101001:ColourData=12'h242;
20'b00000100000000101001:ColourData=12'h0F0;
20'b00000100010000101001:ColourData=12'h2D0;
20'b00000100100000101001:ColourData=12'h4A0;
20'b00000100110000101001:ColourData=12'hA40;
20'b00000101000000101001:ColourData=12'hA30;
20'b00000101010000101001:ColourData=12'hB40;
20'b00000101100000101001:ColourData=12'hE50;
20'b00000101110000101001:ColourData=12'hE50;
20'b00000110000000101001:ColourData=12'hE50;
20'b00000110010000101001:ColourData=12'hD40;
20'b00000110100000101001:ColourData=12'hA30;
20'b00000110110000101001:ColourData=12'hA30;
20'b00000111000000101001:ColourData=12'h770;
20'b00000111010000101001:ColourData=12'h2C0;
20'b00000111100000101001:ColourData=12'h1E0;
20'b00000111110000101001:ColourData=12'h6F6;
20'b00000000000000101010:ColourData=12'hD99;
20'b00000000010000101010:ColourData=12'hD77;
20'b00000000100000101010:ColourData=12'hD77;
20'b00000000110000101010:ColourData=12'hD77;
20'b00000001000000101010:ColourData=12'h841;
20'b00000001010000101010:ColourData=12'h730;
20'b00000001100000101010:ColourData=12'h730;
20'b00000001110000101010:ColourData=12'h730;
20'b00000010000000101010:ColourData=12'h730;
20'b00000010010000101010:ColourData=12'h730;
20'b00000010100000101010:ColourData=12'h730;
20'b00000010110000101010:ColourData=12'h630;
20'b00000011000000101010:ColourData=12'h000;
20'b00000011010000101010:ColourData=12'h000;
20'b00000011100000101010:ColourData=12'h000;
20'b00000011110000101010:ColourData=12'h242;
20'b00000100000000101010:ColourData=12'h5B1;
20'b00000100010000101010:ColourData=12'hD50;
20'b00000100100000101010:ColourData=12'hB63;
20'b00000100110000101010:ColourData=12'h443;
20'b00000101000000101010:ColourData=12'h444;
20'b00000101010000101010:ColourData=12'h643;
20'b00000101100000101010:ColourData=12'hA40;
20'b00000101110000101010:ColourData=12'hA40;
20'b00000110000000101010:ColourData=12'hA40;
20'b00000110010000101010:ColourData=12'h841;
20'b00000110100000101010:ColourData=12'h443;
20'b00000110110000101010:ColourData=12'h443;
20'b00000111000000101010:ColourData=12'h853;
20'b00000111010000101010:ColourData=12'hE62;
20'b00000111100000101010:ColourData=12'h880;
20'b00000111110000101010:ColourData=12'h7E6;
20'b00000000000000101011:ColourData=12'hD99;
20'b00000000010000101011:ColourData=12'hD77;
20'b00000000100000101011:ColourData=12'hD77;
20'b00000000110000101011:ColourData=12'hB66;
20'b00000001000000101011:ColourData=12'h731;
20'b00000001010000101011:ColourData=12'h630;
20'b00000001100000101011:ColourData=12'h630;
20'b00000001110000101011:ColourData=12'h630;
20'b00000010000000101011:ColourData=12'h630;
20'b00000010010000101011:ColourData=12'h630;
20'b00000010100000101011:ColourData=12'h630;
20'b00000010110000101011:ColourData=12'h520;
20'b00000011000000101011:ColourData=12'h000;
20'b00000011010000101011:ColourData=12'h000;
20'b00000011100000101011:ColourData=12'h000;
20'b00000011110000101011:ColourData=12'h322;
20'b00000100000000101011:ColourData=12'hE51;
20'b00000100010000101011:ColourData=12'hE52;
20'b00000100100000101011:ColourData=12'hEA8;
20'b00000100110000101011:ColourData=12'hEA8;
20'b00000101000000101011:ColourData=12'hEA8;
20'b00000101010000101011:ColourData=12'hB86;
20'b00000101100000101011:ColourData=12'h421;
20'b00000101110000101011:ColourData=12'h420;
20'b00000110000000101011:ColourData=12'h410;
20'b00000110010000101011:ColourData=12'h743;
20'b00000110100000101011:ColourData=12'hEA8;
20'b00000110110000101011:ColourData=12'hEA8;
20'b00000111000000101011:ColourData=12'hEA8;
20'b00000111010000101011:ColourData=12'hE85;
20'b00000111100000101011:ColourData=12'hE40;
20'b00000111110000101011:ColourData=12'hE96;
20'b00000000000000101100:ColourData=12'hD99;
20'b00000000010000101100:ColourData=12'hD77;
20'b00000000100000101100:ColourData=12'hB66;
20'b00000000110000101100:ColourData=12'h211;
20'b00000001000000101100:ColourData=12'h000;
20'b00000001010000101100:ColourData=12'h000;
20'b00000001100000101100:ColourData=12'h000;
20'b00000001110000101100:ColourData=12'h000;
20'b00000010000000101100:ColourData=12'h000;
20'b00000010010000101100:ColourData=12'h000;
20'b00000010100000101100:ColourData=12'h000;
20'b00000010110000101100:ColourData=12'h000;
20'b00000011000000101100:ColourData=12'h420;
20'b00000011010000101100:ColourData=12'h000;
20'b00000011100000101100:ColourData=12'h000;
20'b00000011110000101100:ColourData=12'h332;
20'b00000100000000101100:ColourData=12'hB81;
20'b00000100010000101100:ColourData=12'hA70;
20'b00000100100000101100:ColourData=12'hB71;
20'b00000100110000101100:ColourData=12'hE63;
20'b00000101000000101100:ColourData=12'hE63;
20'b00000101010000101100:ColourData=12'hE62;
20'b00000101100000101100:ColourData=12'hD62;
20'b00000101110000101100:ColourData=12'hD62;
20'b00000110000000101100:ColourData=12'hD62;
20'b00000110010000101100:ColourData=12'hD62;
20'b00000110100000101100:ColourData=12'hE63;
20'b00000110110000101100:ColourData=12'hE63;
20'b00000111000000101100:ColourData=12'hD72;
20'b00000111010000101100:ColourData=12'hA70;
20'b00000111100000101100:ColourData=12'hA70;
20'b00000111110000101100:ColourData=12'hCA6;
20'b00000000000000101101:ColourData=12'hD99;
20'b00000000010000101101:ColourData=12'hB66;
20'b00000000100000101101:ColourData=12'h211;
20'b00000000110000101101:ColourData=12'h000;
20'b00000001000000101101:ColourData=12'h000;
20'b00000001010000101101:ColourData=12'h000;
20'b00000001100000101101:ColourData=12'h000;
20'b00000001110000101101:ColourData=12'h000;
20'b00000010000000101101:ColourData=12'h000;
20'b00000010010000101101:ColourData=12'h000;
20'b00000010100000101101:ColourData=12'h000;
20'b00000010110000101101:ColourData=12'h000;
20'b00000011000000101101:ColourData=12'h000;
20'b00000011010000101101:ColourData=12'h420;
20'b00000011100000101101:ColourData=12'h000;
20'b00000011110000101101:ColourData=12'h242;
20'b00000100000000101101:ColourData=12'h0F0;
20'b00000100010000101101:ColourData=12'h0F0;
20'b00000100100000101101:ColourData=12'h2F1;
20'b00000100110000101101:ColourData=12'hBD8;
20'b00000101000000101101:ColourData=12'hFCA;
20'b00000101010000101101:ColourData=12'hFCA;
20'b00000101100000101101:ColourData=12'hFCA;
20'b00000101110000101101:ColourData=12'hFCA;
20'b00000110000000101101:ColourData=12'hFCA;
20'b00000110010000101101:ColourData=12'hFCA;
20'b00000110100000101101:ColourData=12'hFCA;
20'b00000110110000101101:ColourData=12'hEDA;
20'b00000111000000101101:ColourData=12'h7E4;
20'b00000111010000101101:ColourData=12'h0F0;
20'b00000111100000101101:ColourData=12'h0F0;
20'b00000111110000101101:ColourData=12'h6F6;
20'b00000000000000101110:ColourData=12'hC88;
20'b00000000010000101110:ColourData=12'h311;
20'b00000000100000101110:ColourData=12'h000;
20'b00000000110000101110:ColourData=12'h000;
20'b00000001000000101110:ColourData=12'h000;
20'b00000001010000101110:ColourData=12'h000;
20'b00000001100000101110:ColourData=12'h000;
20'b00000001110000101110:ColourData=12'h000;
20'b00000010000000101110:ColourData=12'h000;
20'b00000010010000101110:ColourData=12'h000;
20'b00000010100000101110:ColourData=12'h000;
20'b00000010110000101110:ColourData=12'h000;
20'b00000011000000101110:ColourData=12'h000;
20'b00000011010000101110:ColourData=12'h000;
20'b00000011100000101110:ColourData=12'h410;
20'b00000011110000101110:ColourData=12'h342;
20'b00000100000000101110:ColourData=12'h0E0;
20'b00000100010000101110:ColourData=12'h0C0;
20'b00000100100000101110:ColourData=12'h0B0;
20'b00000100110000101110:ColourData=12'h2B2;
20'b00000101000000101110:ColourData=12'hBA8;
20'b00000101010000101110:ColourData=12'hBB8;
20'b00000101100000101110:ColourData=12'hAD8;
20'b00000101110000101110:ColourData=12'hAD8;
20'b00000110000000101110:ColourData=12'hAD8;
20'b00000110010000101110:ColourData=12'hBC8;
20'b00000110100000101110:ColourData=12'hC99;
20'b00000110110000101110:ColourData=12'h7A5;
20'b00000111000000101110:ColourData=12'h0B0;
20'b00000111010000101110:ColourData=12'h0B0;
20'b00000111100000101110:ColourData=12'h0D0;
20'b00000111110000101110:ColourData=12'h6F6;
20'b00000000000000101111:ColourData=12'h433;
20'b00000000010000101111:ColourData=12'h000;
20'b00000000100000101111:ColourData=12'h000;
20'b00000000110000101111:ColourData=12'h000;
20'b00000001000000101111:ColourData=12'h000;
20'b00000001010000101111:ColourData=12'h000;
20'b00000001100000101111:ColourData=12'h000;
20'b00000001110000101111:ColourData=12'h000;
20'b00000010000000101111:ColourData=12'h000;
20'b00000010010000101111:ColourData=12'h000;
20'b00000010100000101111:ColourData=12'h000;
20'b00000010110000101111:ColourData=12'h000;
20'b00000011000000101111:ColourData=12'h000;
20'b00000011010000101111:ColourData=12'h000;
20'b00000011100000101111:ColourData=12'h000;
20'b00000011110000101111:ColourData=12'h662;
20'b00000100000000101111:ColourData=12'h0D0;
20'b00000100010000101111:ColourData=12'h050;
20'b00000100100000101111:ColourData=12'h041;
20'b00000100110000101111:ColourData=12'h141;
20'b00000101000000101111:ColourData=12'h411;
20'b00000101010000101111:ColourData=12'h440;
20'b00000101100000101111:ColourData=12'h3C0;
20'b00000101110000101111:ColourData=12'h3C0;
20'b00000110000000101111:ColourData=12'h3C0;
20'b00000110010000101111:ColourData=12'h2A0;
20'b00000110100000101111:ColourData=12'h051;
20'b00000110110000101111:ColourData=12'h051;
20'b00000111000000101111:ColourData=12'h050;
20'b00000111010000101111:ColourData=12'h141;
20'b00000111100000101111:ColourData=12'h080;
20'b00000111110000101111:ColourData=12'h6F6;
20'b00000000000000110000:ColourData=12'h222;
20'b00000000010000110000:ColourData=12'h000;
20'b00000000100000110000:ColourData=12'h010;
20'b00000000110000110000:ColourData=12'h010;
20'b00000001000000110000:ColourData=12'h010;
20'b00000001010000110000:ColourData=12'h010;
20'b00000001100000110000:ColourData=12'h010;
20'b00000001110000110000:ColourData=12'h010;
20'b00000010000000110000:ColourData=12'h010;
20'b00000010010000110000:ColourData=12'h010;
20'b00000010100000110000:ColourData=12'h010;
20'b00000010110000110000:ColourData=12'h010;
20'b00000011000000110000:ColourData=12'h010;
20'b00000011010000110000:ColourData=12'h010;
20'b00000011100000110000:ColourData=12'h010;
20'b00000011110000110000:ColourData=12'h252;
20'b00000100000000110000:ColourData=12'h0F0;
20'b00000100010000110000:ColourData=12'h0F0;
20'b00000100100000110000:ColourData=12'h0E0;
20'b00000100110000110000:ColourData=12'h5A0;
20'b00000101000000110000:ColourData=12'hE20;
20'b00000101010000110000:ColourData=12'hF20;
20'b00000101100000110000:ColourData=12'hE30;
20'b00000101110000110000:ColourData=12'hE20;
20'b00000110000000110000:ColourData=12'hF20;
20'b00000110010000110000:ColourData=12'hB50;
20'b00000110100000110000:ColourData=12'h3C0;
20'b00000110110000110000:ColourData=12'h3B0;
20'b00000111000000110000:ColourData=12'h2D0;
20'b00000111010000110000:ColourData=12'h0F0;
20'b00000111100000110000:ColourData=12'h0F0;
20'b00000111110000110000:ColourData=12'h6F6;
20'b00000000000000110001:ColourData=12'h333;
20'b00000000010000110001:ColourData=12'h290;
20'b00000000100000110001:ColourData=12'h3D1;
20'b00000000110000110001:ColourData=12'h3D1;
20'b00000001000000110001:ColourData=12'h3D1;
20'b00000001010000110001:ColourData=12'h3D1;
20'b00000001100000110001:ColourData=12'h3D1;
20'b00000001110000110001:ColourData=12'h3D1;
20'b00000010000000110001:ColourData=12'h3D1;
20'b00000010010000110001:ColourData=12'h3D1;
20'b00000010100000110001:ColourData=12'h3D1;
20'b00000010110000110001:ColourData=12'h3D1;
20'b00000011000000110001:ColourData=12'h3D1;
20'b00000011010000110001:ColourData=12'h3D1;
20'b00000011100000110001:ColourData=12'h3D1;
20'b00000011110000110001:ColourData=12'h4D3;
20'b00000100000000110001:ColourData=12'h0F0;
20'b00000100010000110001:ColourData=12'h0F0;
20'b00000100100000110001:ColourData=12'h2D0;
20'b00000100110000110001:ColourData=12'hD40;
20'b00000101000000110001:ColourData=12'hD30;
20'b00000101010000110001:ColourData=12'hD30;
20'b00000101100000110001:ColourData=12'hE40;
20'b00000101110000110001:ColourData=12'hF40;
20'b00000110000000110001:ColourData=12'hE40;
20'b00000110010000110001:ColourData=12'hE40;
20'b00000110100000110001:ColourData=12'hD50;
20'b00000110110000110001:ColourData=12'hB50;
20'b00000111000000110001:ColourData=12'h690;
20'b00000111010000110001:ColourData=12'h0F0;
20'b00000111100000110001:ColourData=12'h0F0;
20'b00000111110000110001:ColourData=12'h6F6;
20'b00000000000000110010:ColourData=12'h333;
20'b00000000010000110010:ColourData=12'h160;
20'b00000000100000110010:ColourData=12'h290;
20'b00000000110000110010:ColourData=12'h290;
20'b00000001000000110010:ColourData=12'h280;
20'b00000001010000110010:ColourData=12'h280;
20'b00000001100000110010:ColourData=12'h3E1;
20'b00000001110000110010:ColourData=12'h4F1;
20'b00000010000000110010:ColourData=12'h3F1;
20'b00000010010000110010:ColourData=12'h3F1;
20'b00000010100000110010:ColourData=12'h3F1;
20'b00000010110000110010:ColourData=12'h3F1;
20'b00000011000000110010:ColourData=12'h290;
20'b00000011010000110010:ColourData=12'h290;
20'b00000011100000110010:ColourData=12'h280;
20'b00000011110000110010:ColourData=12'h3A2;
20'b00000100000000110010:ColourData=12'h0F0;
20'b00000100010000110010:ColourData=12'h0F0;
20'b00000100100000110010:ColourData=12'h3C0;
20'b00000100110000110010:ColourData=12'hA70;
20'b00000101000000110010:ColourData=12'hB70;
20'b00000101010000110010:ColourData=12'hA70;
20'b00000101100000110010:ColourData=12'hC81;
20'b00000101110000110010:ColourData=12'hF93;
20'b00000110000000110010:ColourData=12'hD82;
20'b00000110010000110010:ColourData=12'hC70;
20'b00000110100000110010:ColourData=12'hBB2;
20'b00000110110000110010:ColourData=12'h3D0;
20'b00000111000000110010:ColourData=12'h1E0;
20'b00000111010000110010:ColourData=12'h0F0;
20'b00000111100000110010:ColourData=12'h0F0;
20'b00000111110000110010:ColourData=12'h6F6;
20'b00000000000000110011:ColourData=12'h333;
20'b00000000010000110011:ColourData=12'h2A0;
20'b00000000100000110011:ColourData=12'h3E1;
20'b00000000110000110011:ColourData=12'h3E1;
20'b00000001000000110011:ColourData=12'h280;
20'b00000001010000110011:ColourData=12'h170;
20'b00000001100000110011:ColourData=12'h3E1;
20'b00000001110000110011:ColourData=12'h3F1;
20'b00000010000000110011:ColourData=12'h3F1;
20'b00000010010000110011:ColourData=12'h3F1;
20'b00000010100000110011:ColourData=12'h3F1;
20'b00000010110000110011:ColourData=12'h3E1;
20'b00000011000000110011:ColourData=12'h280;
20'b00000011010000110011:ColourData=12'h3D1;
20'b00000011100000110011:ColourData=12'h3D1;
20'b00000011110000110011:ColourData=12'h3A2;
20'b00000100000000110011:ColourData=12'h0F0;
20'b00000100010000110011:ColourData=12'h1D0;
20'b00000100100000110011:ColourData=12'h970;
20'b00000100110000110011:ColourData=12'hB70;
20'b00000101000000110011:ColourData=12'hE92;
20'b00000101010000110011:ColourData=12'hB70;
20'b00000101100000110011:ColourData=12'hE92;
20'b00000101110000110011:ColourData=12'hF93;
20'b00000110000000110011:ColourData=12'hE92;
20'b00000110010000110011:ColourData=12'hC81;
20'b00000110100000110011:ColourData=12'hE92;
20'b00000110110000110011:ColourData=12'hF93;
20'b00000111000000110011:ColourData=12'hBB2;
20'b00000111010000110011:ColourData=12'h2E0;
20'b00000111100000110011:ColourData=12'h0F0;
20'b00000111110000110011:ColourData=12'h6F6;
20'b00000000000000110100:ColourData=12'h333;
20'b00000000010000110100:ColourData=12'h2B0;
20'b00000000100000110100:ColourData=12'h4F1;
20'b00000000110000110100:ColourData=12'h3F1;
20'b00000001000000110100:ColourData=12'h280;
20'b00000001010000110100:ColourData=12'h170;
20'b00000001100000110100:ColourData=12'h3E1;
20'b00000001110000110100:ColourData=12'h3F1;
20'b00000010000000110100:ColourData=12'h3F1;
20'b00000010010000110100:ColourData=12'h3F1;
20'b00000010100000110100:ColourData=12'h3F1;
20'b00000010110000110100:ColourData=12'h3E1;
20'b00000011000000110100:ColourData=12'h290;
20'b00000011010000110100:ColourData=12'h3E1;
20'b00000011100000110100:ColourData=12'h3E1;
20'b00000011110000110100:ColourData=12'h3A2;
20'b00000100000000110100:ColourData=12'h0F0;
20'b00000100010000110100:ColourData=12'h1D0;
20'b00000100100000110100:ColourData=12'hA70;
20'b00000100110000110100:ColourData=12'hB70;
20'b00000101000000110100:ColourData=12'hD81;
20'b00000101010000110100:ColourData=12'hB70;
20'b00000101100000110100:ColourData=12'hC81;
20'b00000101110000110100:ColourData=12'hF93;
20'b00000110000000110100:ColourData=12'hF93;
20'b00000110010000110100:ColourData=12'hC81;
20'b00000110100000110100:ColourData=12'hB70;
20'b00000110110000110100:ColourData=12'hE92;
20'b00000111000000110100:ColourData=12'hD92;
20'b00000111010000110100:ColourData=12'h7C1;
20'b00000111100000110100:ColourData=12'h0F0;
20'b00000111110000110100:ColourData=12'h6F6;
20'b00000000000000110101:ColourData=12'h333;
20'b00000000010000110101:ColourData=12'h2B0;
20'b00000000100000110101:ColourData=12'h4F1;
20'b00000000110000110101:ColourData=12'h3F1;
20'b00000001000000110101:ColourData=12'h280;
20'b00000001010000110101:ColourData=12'h170;
20'b00000001100000110101:ColourData=12'h3E1;
20'b00000001110000110101:ColourData=12'h3F1;
20'b00000010000000110101:ColourData=12'h3F1;
20'b00000010010000110101:ColourData=12'h3F1;
20'b00000010100000110101:ColourData=12'h3F1;
20'b00000010110000110101:ColourData=12'h3E1;
20'b00000011000000110101:ColourData=12'h290;
20'b00000011010000110101:ColourData=12'h3E1;
20'b00000011100000110101:ColourData=12'h3E1;
20'b00000011110000110101:ColourData=12'h3A2;
20'b00000100000000110101:ColourData=12'h0F0;
20'b00000100010000110101:ColourData=12'h1E0;
20'b00000100100000110101:ColourData=12'h790;
20'b00000100110000110101:ColourData=12'h880;
20'b00000101000000110101:ColourData=12'hC81;
20'b00000101010000110101:ColourData=12'hF93;
20'b00000101100000110101:ColourData=12'hF93;
20'b00000101110000110101:ColourData=12'hF93;
20'b00000110000000110101:ColourData=12'hE92;
20'b00000110010000110101:ColourData=12'hB70;
20'b00000110100000110101:ColourData=12'hB70;
20'b00000110110000110101:ColourData=12'hA70;
20'b00000111000000110101:ColourData=12'h4B0;
20'b00000111010000110101:ColourData=12'h0F0;
20'b00000111100000110101:ColourData=12'h0F0;
20'b00000111110000110101:ColourData=12'h6F6;
20'b00000000000000110110:ColourData=12'h333;
20'b00000000010000110110:ColourData=12'h2B0;
20'b00000000100000110110:ColourData=12'h4F1;
20'b00000000110000110110:ColourData=12'h3F1;
20'b00000001000000110110:ColourData=12'h280;
20'b00000001010000110110:ColourData=12'h170;
20'b00000001100000110110:ColourData=12'h3E1;
20'b00000001110000110110:ColourData=12'h3F1;
20'b00000010000000110110:ColourData=12'h3F1;
20'b00000010010000110110:ColourData=12'h3F1;
20'b00000010100000110110:ColourData=12'h3F1;
20'b00000010110000110110:ColourData=12'h3E1;
20'b00000011000000110110:ColourData=12'h290;
20'b00000011010000110110:ColourData=12'h3E1;
20'b00000011100000110110:ColourData=12'h3E1;
20'b00000011110000110110:ColourData=12'h3A2;
20'b00000100000000110110:ColourData=12'h0F0;
20'b00000100010000110110:ColourData=12'h0F0;
20'b00000100100000110110:ColourData=12'h0F0;
20'b00000100110000110110:ColourData=12'h4C0;
20'b00000101000000110110:ColourData=12'hE92;
20'b00000101010000110110:ColourData=12'hE82;
20'b00000101100000110110:ColourData=12'hF82;
20'b00000101110000110110:ColourData=12'hE92;
20'b00000110000000110110:ColourData=12'hE92;
20'b00000110010000110110:ColourData=12'hD92;
20'b00000110100000110110:ColourData=12'hBB2;
20'b00000110110000110110:ColourData=12'h7C1;
20'b00000111000000110110:ColourData=12'h0F0;
20'b00000111010000110110:ColourData=12'h0F0;
20'b00000111100000110110:ColourData=12'h0F0;
20'b00000111110000110110:ColourData=12'h6F6;
20'b00000000000000110111:ColourData=12'h333;
20'b00000000010000110111:ColourData=12'h2B0;
20'b00000000100000110111:ColourData=12'h4F1;
20'b00000000110000110111:ColourData=12'h3F1;
20'b00000001000000110111:ColourData=12'h280;
20'b00000001010000110111:ColourData=12'h170;
20'b00000001100000110111:ColourData=12'h3E1;
20'b00000001110000110111:ColourData=12'h3F1;
20'b00000010000000110111:ColourData=12'h3F1;
20'b00000010010000110111:ColourData=12'h3F1;
20'b00000010100000110111:ColourData=12'h3F1;
20'b00000010110000110111:ColourData=12'h3E1;
20'b00000011000000110111:ColourData=12'h290;
20'b00000011010000110111:ColourData=12'h3E1;
20'b00000011100000110111:ColourData=12'h3E1;
20'b00000011110000110111:ColourData=12'h3A2;
20'b00000100000000110111:ColourData=12'h0F0;
20'b00000100010000110111:ColourData=12'h0F0;
20'b00000100100000110111:ColourData=12'h3C0;
20'b00000100110000110111:ColourData=12'hA70;
20'b00000101000000110111:ColourData=12'hA70;
20'b00000101010000110111:ColourData=12'hB60;
20'b00000101100000110111:ColourData=12'hD40;
20'b00000101110000110111:ColourData=12'hA70;
20'b00000110000000110111:ColourData=12'hA60;
20'b00000110010000110111:ColourData=12'h880;
20'b00000110100000110111:ColourData=12'h2D0;
20'b00000110110000110111:ColourData=12'h2D0;
20'b00000111000000110111:ColourData=12'h0E0;
20'b00000111010000110111:ColourData=12'h0F0;
20'b00000111100000110111:ColourData=12'h0F0;
20'b00000111110000110111:ColourData=12'h6F6;
20'b00000000000000111000:ColourData=12'h333;
20'b00000000010000111000:ColourData=12'h2B0;
20'b00000000100000111000:ColourData=12'h4F1;
20'b00000000110000111000:ColourData=12'h3F1;
20'b00000001000000111000:ColourData=12'h280;
20'b00000001010000111000:ColourData=12'h170;
20'b00000001100000111000:ColourData=12'h3E1;
20'b00000001110000111000:ColourData=12'h3F1;
20'b00000010000000111000:ColourData=12'h3F1;
20'b00000010010000111000:ColourData=12'h3F1;
20'b00000010100000111000:ColourData=12'h3F1;
20'b00000010110000111000:ColourData=12'h3E1;
20'b00000011000000111000:ColourData=12'h290;
20'b00000011010000111000:ColourData=12'h3E1;
20'b00000011100000111000:ColourData=12'h3E1;
20'b00000011110000111000:ColourData=12'h3A2;
20'b00000100000000111000:ColourData=12'h0F0;
20'b00000100010000111000:ColourData=12'h3C0;
20'b00000100100000111000:ColourData=12'h970;
20'b00000100110000111000:ColourData=12'hA70;
20'b00000101000000111000:ColourData=12'hA70;
20'b00000101010000111000:ColourData=12'hB60;
20'b00000101100000111000:ColourData=12'hE30;
20'b00000101110000111000:ColourData=12'hB60;
20'b00000110000000111000:ColourData=12'hC50;
20'b00000110010000111000:ColourData=12'hD40;
20'b00000110100000111000:ColourData=12'h970;
20'b00000110110000111000:ColourData=12'hA70;
20'b00000111000000111000:ColourData=12'h790;
20'b00000111010000111000:ColourData=12'h0E0;
20'b00000111100000111000:ColourData=12'h0F0;
20'b00000111110000111000:ColourData=12'h6F6;
20'b00000000000000111001:ColourData=12'h333;
20'b00000000010000111001:ColourData=12'h2B0;
20'b00000000100000111001:ColourData=12'h4F1;
20'b00000000110000111001:ColourData=12'h3F1;
20'b00000001000000111001:ColourData=12'h280;
20'b00000001010000111001:ColourData=12'h170;
20'b00000001100000111001:ColourData=12'h3E1;
20'b00000001110000111001:ColourData=12'h3F1;
20'b00000010000000111001:ColourData=12'h3F1;
20'b00000010010000111001:ColourData=12'h3F1;
20'b00000010100000111001:ColourData=12'h3F1;
20'b00000010110000111001:ColourData=12'h3E1;
20'b00000011000000111001:ColourData=12'h290;
20'b00000011010000111001:ColourData=12'h3E1;
20'b00000011100000111001:ColourData=12'h3E1;
20'b00000011110000111001:ColourData=12'h3A2;
20'b00000100000000111001:ColourData=12'h2E0;
20'b00000100010000111001:ColourData=12'hB80;
20'b00000100100000111001:ColourData=12'hB70;
20'b00000100110000111001:ColourData=12'hB70;
20'b00000101000000111001:ColourData=12'hA70;
20'b00000101010000111001:ColourData=12'hC50;
20'b00000101100000111001:ColourData=12'hF40;
20'b00000101110000111001:ColourData=12'hE20;
20'b00000110000000111001:ColourData=12'hF30;
20'b00000110010000111001:ColourData=12'hE50;
20'b00000110100000111001:ColourData=12'hA60;
20'b00000110110000111001:ColourData=12'hA70;
20'b00000111000000111001:ColourData=12'hB70;
20'b00000111010000111001:ColourData=12'h6A0;
20'b00000111100000111001:ColourData=12'h0F0;
20'b00000111110000111001:ColourData=12'h6F6;
20'b00000000000000111010:ColourData=12'h333;
20'b00000000010000111010:ColourData=12'h2B0;
20'b00000000100000111010:ColourData=12'h4F1;
20'b00000000110000111010:ColourData=12'h3F1;
20'b00000001000000111010:ColourData=12'h280;
20'b00000001010000111010:ColourData=12'h170;
20'b00000001100000111010:ColourData=12'h3E1;
20'b00000001110000111010:ColourData=12'h3F1;
20'b00000010000000111010:ColourData=12'h3F1;
20'b00000010010000111010:ColourData=12'h3F1;
20'b00000010100000111010:ColourData=12'h3F1;
20'b00000010110000111010:ColourData=12'h3E1;
20'b00000011000000111010:ColourData=12'h290;
20'b00000011010000111010:ColourData=12'h3E1;
20'b00000011100000111010:ColourData=12'h3E1;
20'b00000011110000111010:ColourData=12'h3A2;
20'b00000100000000111010:ColourData=12'h3E1;
20'b00000100010000111010:ColourData=12'hE93;
20'b00000100100000111010:ColourData=12'hF93;
20'b00000100110000111010:ColourData=12'hE92;
20'b00000101000000111010:ColourData=12'hC60;
20'b00000101010000111010:ColourData=12'hF40;
20'b00000101100000111010:ColourData=12'hF61;
20'b00000101110000111010:ColourData=12'hF20;
20'b00000110000000111010:ColourData=12'hF40;
20'b00000110010000111010:ColourData=12'hF61;
20'b00000110100000111010:ColourData=12'hD40;
20'b00000110110000111010:ColourData=12'hC81;
20'b00000111000000111010:ColourData=12'hF93;
20'b00000111010000111010:ColourData=12'h9B2;
20'b00000111100000111010:ColourData=12'h0F0;
20'b00000111110000111010:ColourData=12'h6F6;
20'b00000000000000111011:ColourData=12'h333;
20'b00000000010000111011:ColourData=12'h2B0;
20'b00000000100000111011:ColourData=12'h4F1;
20'b00000000110000111011:ColourData=12'h3F1;
20'b00000001000000111011:ColourData=12'h280;
20'b00000001010000111011:ColourData=12'h170;
20'b00000001100000111011:ColourData=12'h3E1;
20'b00000001110000111011:ColourData=12'h3F1;
20'b00000010000000111011:ColourData=12'h3F1;
20'b00000010010000111011:ColourData=12'h3F1;
20'b00000010100000111011:ColourData=12'h3F1;
20'b00000010110000111011:ColourData=12'h3E1;
20'b00000011000000111011:ColourData=12'h290;
20'b00000011010000111011:ColourData=12'h3E1;
20'b00000011100000111011:ColourData=12'h3E1;
20'b00000011110000111011:ColourData=12'h3A2;
20'b00000100000000111011:ColourData=12'h3E1;
20'b00000100010000111011:ColourData=12'hF93;
20'b00000100100000111011:ColourData=12'hF93;
20'b00000100110000111011:ColourData=12'hF93;
20'b00000101000000111011:ColourData=12'hF61;
20'b00000101010000111011:ColourData=12'hF30;
20'b00000101100000111011:ColourData=12'hF20;
20'b00000101110000111011:ColourData=12'hF20;
20'b00000110000000111011:ColourData=12'hF30;
20'b00000110010000111011:ColourData=12'hF20;
20'b00000110100000111011:ColourData=12'hF40;
20'b00000110110000111011:ColourData=12'hF82;
20'b00000111000000111011:ColourData=12'hF93;
20'b00000111010000111011:ColourData=12'h9B2;
20'b00000111100000111011:ColourData=12'h0F0;
20'b00000111110000111011:ColourData=12'h6F6;
20'b00000000000000111100:ColourData=12'h333;
20'b00000000010000111100:ColourData=12'h2B0;
20'b00000000100000111100:ColourData=12'h4F1;
20'b00000000110000111100:ColourData=12'h3F1;
20'b00000001000000111100:ColourData=12'h290;
20'b00000001010000111100:ColourData=12'h170;
20'b00000001100000111100:ColourData=12'h3E1;
20'b00000001110000111100:ColourData=12'h4F1;
20'b00000010000000111100:ColourData=12'h3F1;
20'b00000010010000111100:ColourData=12'h3F1;
20'b00000010100000111100:ColourData=12'h3F1;
20'b00000010110000111100:ColourData=12'h3E1;
20'b00000011000000111100:ColourData=12'h290;
20'b00000011010000111100:ColourData=12'h3E1;
20'b00000011100000111100:ColourData=12'h3E1;
20'b00000011110000111100:ColourData=12'h3A2;
20'b00000100000000111100:ColourData=12'h2E0;
20'b00000100010000111100:ColourData=12'hBB2;
20'b00000100100000111100:ColourData=12'hCA2;
20'b00000100110000111100:ColourData=12'hF61;
20'b00000101000000111100:ColourData=12'hF30;
20'b00000101010000111100:ColourData=12'hF20;
20'b00000101100000111100:ColourData=12'hE30;
20'b00000101110000111100:ColourData=12'hC40;
20'b00000110000000111100:ColourData=12'hF20;
20'b00000110010000111100:ColourData=12'hF20;
20'b00000110100000111100:ColourData=12'hF20;
20'b00000110110000111100:ColourData=12'hD50;
20'b00000111000000111100:ColourData=12'hBB2;
20'b00000111010000111100:ColourData=12'h7C1;
20'b00000111100000111100:ColourData=12'h0F0;
20'b00000111110000111100:ColourData=12'h6F6;
20'b00000000000000111101:ColourData=12'h323;
20'b00000000010000111101:ColourData=12'h2A0;
20'b00000000100000111101:ColourData=12'h3D1;
20'b00000000110000111101:ColourData=12'h3D1;
20'b00000001000000111101:ColourData=12'h180;
20'b00000001010000111101:ColourData=12'h160;
20'b00000001100000111101:ColourData=12'h3C1;
20'b00000001110000111101:ColourData=12'h3D1;
20'b00000010000000111101:ColourData=12'h3D1;
20'b00000010010000111101:ColourData=12'h3D1;
20'b00000010100000111101:ColourData=12'h3D1;
20'b00000010110000111101:ColourData=12'h3D1;
20'b00000011000000111101:ColourData=12'h180;
20'b00000011010000111101:ColourData=12'h3D1;
20'b00000011100000111101:ColourData=12'h3C1;
20'b00000011110000111101:ColourData=12'h392;
20'b00000100000000111101:ColourData=12'h0F0;
20'b00000100010000111101:ColourData=12'h0F0;
20'b00000100100000111101:ColourData=12'h4B0;
20'b00000100110000111101:ColourData=12'hD40;
20'b00000101000000111101:ColourData=12'hE30;
20'b00000101010000111101:ColourData=12'hD40;
20'b00000101100000111101:ColourData=12'h780;
20'b00000101110000111101:ColourData=12'h2C0;
20'b00000110000000111101:ColourData=12'hC50;
20'b00000110010000111101:ColourData=12'hE30;
20'b00000110100000111101:ColourData=12'hE30;
20'b00000110110000111101:ColourData=12'hA70;
20'b00000111000000111101:ColourData=12'h1E0;
20'b00000111010000111101:ColourData=12'h0F0;
20'b00000111100000111101:ColourData=12'h0F0;
20'b00000111110000111101:ColourData=12'h6F6;
20'b00000000000000111110:ColourData=12'h343;
20'b00000000010000111110:ColourData=12'h020;
20'b00000000100000111110:ColourData=12'h010;
20'b00000000110000111110:ColourData=12'h010;
20'b00000001000000111110:ColourData=12'h000;
20'b00000001010000111110:ColourData=12'h000;
20'b00000001100000111110:ColourData=12'h000;
20'b00000001110000111110:ColourData=12'h010;
20'b00000010000000111110:ColourData=12'h010;
20'b00000010010000111110:ColourData=12'h010;
20'b00000010100000111110:ColourData=12'h010;
20'b00000010110000111110:ColourData=12'h000;
20'b00000011000000111110:ColourData=12'h000;
20'b00000011010000111110:ColourData=12'h000;
20'b00000011100000111110:ColourData=12'h000;
20'b00000011110000111110:ColourData=12'h242;
20'b00000100000000111110:ColourData=12'h0F0;
20'b00000100010000111110:ColourData=12'h3C0;
20'b00000100100000111110:ColourData=12'hA70;
20'b00000100110000111110:ColourData=12'hA60;
20'b00000101000000111110:ColourData=12'hA60;
20'b00000101010000111110:ColourData=12'h790;
20'b00000101100000111110:ColourData=12'h0F0;
20'b00000101110000111110:ColourData=12'h0F0;
20'b00000110000000111110:ColourData=12'h2C0;
20'b00000110010000111110:ColourData=12'hA60;
20'b00000110100000111110:ColourData=12'hA70;
20'b00000110110000111110:ColourData=12'hA60;
20'b00000111000000111110:ColourData=12'h790;
20'b00000111010000111110:ColourData=12'h1E0;
20'b00000111100000111110:ColourData=12'h0F0;
20'b00000111110000111110:ColourData=12'h6F6;
20'b00000000000000111111:ColourData=12'h2C3;
20'b00000000010000111111:ColourData=12'h0B0;
20'b00000000100000111111:ColourData=12'h010;
20'b00000000110000111111:ColourData=12'h000;
20'b00000001000000111111:ColourData=12'h000;
20'b00000001010000111111:ColourData=12'h000;
20'b00000001100000111111:ColourData=12'h000;
20'b00000001110000111111:ColourData=12'h000;
20'b00000010000000111111:ColourData=12'h000;
20'b00000010010000111111:ColourData=12'h000;
20'b00000010100000111111:ColourData=12'h000;
20'b00000010110000111111:ColourData=12'h000;
20'b00000011000000111111:ColourData=12'h000;
20'b00000011010000111111:ColourData=12'h000;
20'b00000011100000111111:ColourData=12'h000;
20'b00000011110000111111:ColourData=12'h142;
20'b00000100000000111111:ColourData=12'h2E0;
20'b00000100010000111111:ColourData=12'h790;
20'b00000100100000111111:ColourData=12'h790;
20'b00000100110000111111:ColourData=12'h790;
20'b00000101000000111111:ColourData=12'h790;
20'b00000101010000111111:ColourData=12'h5B0;
20'b00000101100000111111:ColourData=12'h0F0;
20'b00000101110000111111:ColourData=12'h0F0;
20'b00000110000000111111:ColourData=12'h1D0;
20'b00000110010000111111:ColourData=12'h790;
20'b00000110100000111111:ColourData=12'h790;
20'b00000110110000111111:ColourData=12'h790;
20'b00000111000000111111:ColourData=12'h880;
20'b00000111010000111111:ColourData=12'h4B0;
20'b00000111100000111111:ColourData=12'h0F0;
20'b00000111110000111111:ColourData=12'h6F6;
20'b00000000000001000000:ColourData=12'h353;
20'b00000000010001000000:ColourData=12'h020;
20'b00000000100001000000:ColourData=12'h010;
20'b00000000110001000000:ColourData=12'h010;
20'b00000001000001000000:ColourData=12'h010;
20'b00000001010001000000:ColourData=12'h010;
20'b00000001100001000000:ColourData=12'h010;
20'b00000001110001000000:ColourData=12'h010;
20'b00000010000001000000:ColourData=12'h010;
20'b00000010010001000000:ColourData=12'h010;
20'b00000010100001000000:ColourData=12'h010;
20'b00000010110001000000:ColourData=12'h010;
20'b00000011000001000000:ColourData=12'h010;
20'b00000011010001000000:ColourData=12'h010;
20'b00000011100001000000:ColourData=12'h000;
20'b00000011110001000000:ColourData=12'h242;
20'b00000100000001000000:ColourData=12'h0F0;
20'b00000100010001000000:ColourData=12'h0F0;
20'b00000100100001000000:ColourData=12'h0F0;
20'b00000100110001000000:ColourData=12'h0F0;
20'b00000101000001000000:ColourData=12'h0E0;
20'b00000101010001000000:ColourData=12'h3C0;
20'b00000101100001000000:ColourData=12'h3C0;
20'b00000101110001000000:ColourData=12'h3C0;
20'b00000110000001000000:ColourData=12'h3C0;
20'b00000110010001000000:ColourData=12'h3C0;
20'b00000110100001000000:ColourData=12'h1D0;
20'b00000110110001000000:ColourData=12'h0F0;
20'b00000111000001000000:ColourData=12'h0F0;
20'b00000111010001000000:ColourData=12'h0F0;
20'b00000111100001000000:ColourData=12'h0F0;
20'b00000111110001000000:ColourData=12'h6F6;
20'b00000000000001000001:ColourData=12'h5D4;
20'b00000000010001000001:ColourData=12'h2C0;
20'b00000000100001000001:ColourData=12'h3D1;
20'b00000000110001000001:ColourData=12'h3D1;
20'b00000001000001000001:ColourData=12'h3D1;
20'b00000001010001000001:ColourData=12'h3D1;
20'b00000001100001000001:ColourData=12'h3D1;
20'b00000001110001000001:ColourData=12'h3D1;
20'b00000010000001000001:ColourData=12'h3D1;
20'b00000010010001000001:ColourData=12'h3D1;
20'b00000010100001000001:ColourData=12'h3D1;
20'b00000010110001000001:ColourData=12'h3D1;
20'b00000011000001000001:ColourData=12'h3D1;
20'b00000011010001000001:ColourData=12'h3D1;
20'b00000011100001000001:ColourData=12'h2A0;
20'b00000011110001000001:ColourData=12'h252;
20'b00000100000001000001:ColourData=12'h0F0;
20'b00000100010001000001:ColourData=12'h0F0;
20'b00000100100001000001:ColourData=12'h0F0;
20'b00000100110001000001:ColourData=12'h0E0;
20'b00000101000001000001:ColourData=12'h5A0;
20'b00000101010001000001:ColourData=12'hE30;
20'b00000101100001000001:ColourData=12'hF20;
20'b00000101110001000001:ColourData=12'hE20;
20'b00000110000001000001:ColourData=12'hE20;
20'b00000110010001000001:ColourData=12'hF20;
20'b00000110100001000001:ColourData=12'hA60;
20'b00000110110001000001:ColourData=12'h3C0;
20'b00000111000001000001:ColourData=12'h3C0;
20'b00000111010001000001:ColourData=12'h2D0;
20'b00000111100001000001:ColourData=12'h0F0;
20'b00000111110001000001:ColourData=12'h6F6;
20'b00000000000001000010:ColourData=12'h4A3;
20'b00000000010001000010:ColourData=12'h180;
20'b00000000100001000010:ColourData=12'h180;
20'b00000000110001000010:ColourData=12'h180;
20'b00000001000001000010:ColourData=12'h180;
20'b00000001010001000010:ColourData=12'h180;
20'b00000001100001000010:ColourData=12'h180;
20'b00000001110001000010:ColourData=12'h180;
20'b00000010000001000010:ColourData=12'h280;
20'b00000010010001000010:ColourData=12'h290;
20'b00000010100001000010:ColourData=12'h280;
20'b00000010110001000010:ColourData=12'h290;
20'b00000011000001000010:ColourData=12'h280;
20'b00000011010001000010:ColourData=12'h290;
20'b00000011100001000010:ColourData=12'h170;
20'b00000011110001000010:ColourData=12'h242;
20'b00000100000001000010:ColourData=12'h0F0;
20'b00000100010001000010:ColourData=12'h0F0;
20'b00000100100001000010:ColourData=12'h0F0;
20'b00000100110001000010:ColourData=12'h2D0;
20'b00000101000001000010:ColourData=12'hD40;
20'b00000101010001000010:ColourData=12'hD30;
20'b00000101100001000010:ColourData=12'hE40;
20'b00000101110001000010:ColourData=12'hF40;
20'b00000110000001000010:ColourData=12'hE40;
20'b00000110010001000010:ColourData=12'hE40;
20'b00000110100001000010:ColourData=12'hF40;
20'b00000110110001000010:ColourData=12'hD50;
20'b00000111000001000010:ColourData=12'hB50;
20'b00000111010001000010:ColourData=12'h690;
20'b00000111100001000010:ColourData=12'h0F0;
20'b00000111110001000010:ColourData=12'h6F6;
20'b00000000000001000011:ColourData=12'h493;
20'b00000000010001000011:ColourData=12'h170;
20'b00000000100001000011:ColourData=12'h170;
20'b00000000110001000011:ColourData=12'h170;
20'b00000001000001000011:ColourData=12'h170;
20'b00000001010001000011:ColourData=12'h170;
20'b00000001100001000011:ColourData=12'h170;
20'b00000001110001000011:ColourData=12'h170;
20'b00000010000001000011:ColourData=12'h170;
20'b00000010010001000011:ColourData=12'h3C1;
20'b00000010100001000011:ColourData=12'h290;
20'b00000010110001000011:ColourData=12'h3C1;
20'b00000011000001000011:ColourData=12'h290;
20'b00000011010001000011:ColourData=12'h3E1;
20'b00000011100001000011:ColourData=12'h2C0;
20'b00000011110001000011:ColourData=12'h252;
20'b00000100000001000011:ColourData=12'h0F0;
20'b00000100010001000011:ColourData=12'h0F0;
20'b00000100100001000011:ColourData=12'h0F0;
20'b00000100110001000011:ColourData=12'h4C0;
20'b00000101000001000011:ColourData=12'hB70;
20'b00000101010001000011:ColourData=12'hA70;
20'b00000101100001000011:ColourData=12'hC81;
20'b00000101110001000011:ColourData=12'hF93;
20'b00000110000001000011:ColourData=12'hD82;
20'b00000110010001000011:ColourData=12'hB70;
20'b00000110100001000011:ColourData=12'hF93;
20'b00000110110001000011:ColourData=12'hBB2;
20'b00000111000001000011:ColourData=12'h3D0;
20'b00000111010001000011:ColourData=12'h1E0;
20'b00000111100001000011:ColourData=12'h0F0;
20'b00000111110001000011:ColourData=12'h6F6;
20'b00000000000001000100:ColourData=12'h493;
20'b00000000010001000100:ColourData=12'h170;
20'b00000000100001000100:ColourData=12'h170;
20'b00000000110001000100:ColourData=12'h170;
20'b00000001000001000100:ColourData=12'h170;
20'b00000001010001000100:ColourData=12'h170;
20'b00000001100001000100:ColourData=12'h170;
20'b00000001110001000100:ColourData=12'h170;
20'b00000010000001000100:ColourData=12'h170;
20'b00000010010001000100:ColourData=12'h290;
20'b00000010100001000100:ColourData=12'h3C1;
20'b00000010110001000100:ColourData=12'h2A0;
20'b00000011000001000100:ColourData=12'h3D1;
20'b00000011010001000100:ColourData=12'h3F1;
20'b00000011100001000100:ColourData=12'h3D1;
20'b00000011110001000100:ColourData=12'h252;
20'b00000100000001000100:ColourData=12'h0F0;
20'b00000100010001000100:ColourData=12'h0F0;
20'b00000100100001000100:ColourData=12'h1D0;
20'b00000100110001000100:ColourData=12'hB80;
20'b00000101000001000100:ColourData=12'hE92;
20'b00000101010001000100:ColourData=12'hB70;
20'b00000101100001000100:ColourData=12'hE92;
20'b00000101110001000100:ColourData=12'hF93;
20'b00000110000001000100:ColourData=12'hE92;
20'b00000110010001000100:ColourData=12'hC81;
20'b00000110100001000100:ColourData=12'hE92;
20'b00000110110001000100:ColourData=12'hF93;
20'b00000111000001000100:ColourData=12'hF93;
20'b00000111010001000100:ColourData=12'hBB2;
20'b00000111100001000100:ColourData=12'h1E0;
20'b00000111110001000100:ColourData=12'h6F6;
20'b00000000000001000101:ColourData=12'h493;
20'b00000000010001000101:ColourData=12'h170;
20'b00000000100001000101:ColourData=12'h170;
20'b00000000110001000101:ColourData=12'h170;
20'b00000001000001000101:ColourData=12'h170;
20'b00000001010001000101:ColourData=12'h170;
20'b00000001100001000101:ColourData=12'h170;
20'b00000001110001000101:ColourData=12'h170;
20'b00000010000001000101:ColourData=12'h180;
20'b00000010010001000101:ColourData=12'h3C1;
20'b00000010100001000101:ColourData=12'h2A0;
20'b00000010110001000101:ColourData=12'h3C1;
20'b00000011000001000101:ColourData=12'h2A0;
20'b00000011010001000101:ColourData=12'h3F1;
20'b00000011100001000101:ColourData=12'h3D1;
20'b00000011110001000101:ColourData=12'h252;
20'b00000100000001000101:ColourData=12'h0F0;
20'b00000100010001000101:ColourData=12'h0F0;
20'b00000100100001000101:ColourData=12'h1D0;
20'b00000100110001000101:ColourData=12'hB70;
20'b00000101000001000101:ColourData=12'hD82;
20'b00000101010001000101:ColourData=12'hB70;
20'b00000101100001000101:ColourData=12'hC81;
20'b00000101110001000101:ColourData=12'hF93;
20'b00000110000001000101:ColourData=12'hF93;
20'b00000110010001000101:ColourData=12'hC81;
20'b00000110100001000101:ColourData=12'hB70;
20'b00000110110001000101:ColourData=12'hE92;
20'b00000111000001000101:ColourData=12'hE82;
20'b00000111010001000101:ColourData=12'hD92;
20'b00000111100001000101:ColourData=12'h6C0;
20'b00000111110001000101:ColourData=12'h6F6;
20'b00000000000001000110:ColourData=12'h493;
20'b00000000010001000110:ColourData=12'h170;
20'b00000000100001000110:ColourData=12'h170;
20'b00000000110001000110:ColourData=12'h170;
20'b00000001000001000110:ColourData=12'h170;
20'b00000001010001000110:ColourData=12'h170;
20'b00000001100001000110:ColourData=12'h170;
20'b00000001110001000110:ColourData=12'h170;
20'b00000010000001000110:ColourData=12'h170;
20'b00000010010001000110:ColourData=12'h290;
20'b00000010100001000110:ColourData=12'h3C1;
20'b00000010110001000110:ColourData=12'h2A0;
20'b00000011000001000110:ColourData=12'h3D1;
20'b00000011010001000110:ColourData=12'h3F1;
20'b00000011100001000110:ColourData=12'h3D1;
20'b00000011110001000110:ColourData=12'h252;
20'b00000100000001000110:ColourData=12'h0F0;
20'b00000100010001000110:ColourData=12'h0F0;
20'b00000100100001000110:ColourData=12'h1E0;
20'b00000100110001000110:ColourData=12'h790;
20'b00000101000001000110:ColourData=12'h990;
20'b00000101010001000110:ColourData=12'hF93;
20'b00000101100001000110:ColourData=12'hF93;
20'b00000101110001000110:ColourData=12'hF93;
20'b00000110000001000110:ColourData=12'hE92;
20'b00000110010001000110:ColourData=12'hB70;
20'b00000110100001000110:ColourData=12'hB70;
20'b00000110110001000110:ColourData=12'hB70;
20'b00000111000001000110:ColourData=12'hA80;
20'b00000111010001000110:ColourData=12'h4B0;
20'b00000111100001000110:ColourData=12'h0F0;
20'b00000111110001000110:ColourData=12'h6F6;
20'b00000000000001000111:ColourData=12'h493;
20'b00000000010001000111:ColourData=12'h170;
20'b00000000100001000111:ColourData=12'h170;
20'b00000000110001000111:ColourData=12'h170;
20'b00000001000001000111:ColourData=12'h170;
20'b00000001010001000111:ColourData=12'h170;
20'b00000001100001000111:ColourData=12'h170;
20'b00000001110001000111:ColourData=12'h170;
20'b00000010000001000111:ColourData=12'h180;
20'b00000010010001000111:ColourData=12'h3C1;
20'b00000010100001000111:ColourData=12'h2A0;
20'b00000010110001000111:ColourData=12'h3C1;
20'b00000011000001000111:ColourData=12'h2A0;
20'b00000011010001000111:ColourData=12'h3F1;
20'b00000011100001000111:ColourData=12'h3D1;
20'b00000011110001000111:ColourData=12'h252;
20'b00000100000001000111:ColourData=12'h0F0;
20'b00000100010001000111:ColourData=12'h0F0;
20'b00000100100001000111:ColourData=12'h0F0;
20'b00000100110001000111:ColourData=12'h0F0;
20'b00000101000001000111:ColourData=12'h5C0;
20'b00000101010001000111:ColourData=12'hE92;
20'b00000101100001000111:ColourData=12'hE92;
20'b00000101110001000111:ColourData=12'hE82;
20'b00000110000001000111:ColourData=12'hF82;
20'b00000110010001000111:ColourData=12'hE92;
20'b00000110100001000111:ColourData=12'hE92;
20'b00000110110001000111:ColourData=12'hF93;
20'b00000111000001000111:ColourData=12'h9B2;
20'b00000111010001000111:ColourData=12'h0F0;
20'b00000111100001000111:ColourData=12'h0F0;
20'b00000111110001000111:ColourData=12'h6F6;
20'b00000000000001001000:ColourData=12'h493;
20'b00000000010001001000:ColourData=12'h170;
20'b00000000100001001000:ColourData=12'h170;
20'b00000000110001001000:ColourData=12'h170;
20'b00000001000001001000:ColourData=12'h170;
20'b00000001010001001000:ColourData=12'h170;
20'b00000001100001001000:ColourData=12'h170;
20'b00000001110001001000:ColourData=12'h170;
20'b00000010000001001000:ColourData=12'h170;
20'b00000010010001001000:ColourData=12'h290;
20'b00000010100001001000:ColourData=12'h3C1;
20'b00000010110001001000:ColourData=12'h2A0;
20'b00000011000001001000:ColourData=12'h3D1;
20'b00000011010001001000:ColourData=12'h3F1;
20'b00000011100001001000:ColourData=12'h3D1;
20'b00000011110001001000:ColourData=12'h252;
20'b00000100000001001000:ColourData=12'h0F0;
20'b00000100010001001000:ColourData=12'h0F0;
20'b00000100100001001000:ColourData=12'h0F0;
20'b00000100110001001000:ColourData=12'h4C0;
20'b00000101000001001000:ColourData=12'hA70;
20'b00000101010001001000:ColourData=12'hA70;
20'b00000101100001001000:ColourData=12'hA70;
20'b00000101110001001000:ColourData=12'hB60;
20'b00000110000001001000:ColourData=12'hC40;
20'b00000110010001001000:ColourData=12'hA70;
20'b00000110100001001000:ColourData=12'hC81;
20'b00000110110001001000:ColourData=12'hF93;
20'b00000111000001001000:ColourData=12'hBB2;
20'b00000111010001001000:ColourData=12'h2E0;
20'b00000111100001001000:ColourData=12'h0F0;
20'b00000111110001001000:ColourData=12'h6F6;
20'b00000000000001001001:ColourData=12'h493;
20'b00000000010001001001:ColourData=12'h170;
20'b00000000100001001001:ColourData=12'h170;
20'b00000000110001001001:ColourData=12'h170;
20'b00000001000001001001:ColourData=12'h170;
20'b00000001010001001001:ColourData=12'h170;
20'b00000001100001001001:ColourData=12'h170;
20'b00000001110001001001:ColourData=12'h170;
20'b00000010000001001001:ColourData=12'h180;
20'b00000010010001001001:ColourData=12'h3C1;
20'b00000010100001001001:ColourData=12'h2A0;
20'b00000010110001001001:ColourData=12'h3C1;
20'b00000011000001001001:ColourData=12'h2A0;
20'b00000011010001001001:ColourData=12'h3F1;
20'b00000011100001001001:ColourData=12'h3D1;
20'b00000011110001001001:ColourData=12'h252;
20'b00000100000001001001:ColourData=12'h0F0;
20'b00000100010001001001:ColourData=12'h0F0;
20'b00000100100001001001:ColourData=12'h6D1;
20'b00000100110001001001:ColourData=12'hE92;
20'b00000101000001001001:ColourData=12'hB60;
20'b00000101010001001001:ColourData=12'hA70;
20'b00000101100001001001:ColourData=12'hA70;
20'b00000101110001001001:ColourData=12'hA70;
20'b00000110000001001001:ColourData=12'h970;
20'b00000110010001001001:ColourData=12'hB80;
20'b00000110100001001001:ColourData=12'hFA3;
20'b00000110110001001001:ColourData=12'hF93;
20'b00000111000001001001:ColourData=12'hEA3;
20'b00000111010001001001:ColourData=12'h7C1;
20'b00000111100001001001:ColourData=12'h0F0;
20'b00000111110001001001:ColourData=12'h6F6;
20'b00000000000001001010:ColourData=12'h493;
20'b00000000010001001010:ColourData=12'h170;
20'b00000000100001001010:ColourData=12'h170;
20'b00000000110001001010:ColourData=12'h170;
20'b00000001000001001010:ColourData=12'h170;
20'b00000001010001001010:ColourData=12'h170;
20'b00000001100001001010:ColourData=12'h170;
20'b00000001110001001010:ColourData=12'h170;
20'b00000010000001001010:ColourData=12'h170;
20'b00000010010001001010:ColourData=12'h290;
20'b00000010100001001010:ColourData=12'h3C1;
20'b00000010110001001010:ColourData=12'h2A0;
20'b00000011000001001010:ColourData=12'h3D1;
20'b00000011010001001010:ColourData=12'h3F1;
20'b00000011100001001010:ColourData=12'h3D1;
20'b00000011110001001010:ColourData=12'h252;
20'b00000100000001001010:ColourData=12'h0F0;
20'b00000100010001001010:ColourData=12'h2E0;
20'b00000100100001001010:ColourData=12'hD92;
20'b00000100110001001010:ColourData=12'hE71;
20'b00000101000001001010:ColourData=12'hE30;
20'b00000101010001001010:ColourData=12'hB60;
20'b00000101100001001010:ColourData=12'hB60;
20'b00000101110001001010:ColourData=12'hB60;
20'b00000110000001001010:ColourData=12'hB60;
20'b00000110010001001010:ColourData=12'hC60;
20'b00000110100001001010:ColourData=12'hF82;
20'b00000110110001001010:ColourData=12'hE92;
20'b00000111000001001010:ColourData=12'h7C1;
20'b00000111010001001010:ColourData=12'h0F0;
20'b00000111100001001010:ColourData=12'h0F0;
20'b00000111110001001010:ColourData=12'h6F6;
20'b00000000000001001011:ColourData=12'h493;
20'b00000000010001001011:ColourData=12'h170;
20'b00000000100001001011:ColourData=12'h170;
20'b00000000110001001011:ColourData=12'h170;
20'b00000001000001001011:ColourData=12'h170;
20'b00000001010001001011:ColourData=12'h170;
20'b00000001100001001011:ColourData=12'h170;
20'b00000001110001001011:ColourData=12'h170;
20'b00000010000001001011:ColourData=12'h180;
20'b00000010010001001011:ColourData=12'h3C1;
20'b00000010100001001011:ColourData=12'h2A0;
20'b00000010110001001011:ColourData=12'h3C1;
20'b00000011000001001011:ColourData=12'h2A0;
20'b00000011010001001011:ColourData=12'h3F1;
20'b00000011100001001011:ColourData=12'h3D1;
20'b00000011110001001011:ColourData=12'h252;
20'b00000100000001001011:ColourData=12'h0F0;
20'b00000100010001001011:ColourData=12'h1D0;
20'b00000100100001001011:ColourData=12'hA70;
20'b00000100110001001011:ColourData=12'hC50;
20'b00000101000001001011:ColourData=12'hF30;
20'b00000101010001001011:ColourData=12'hE30;
20'b00000101100001001011:ColourData=12'hE30;
20'b00000101110001001011:ColourData=12'hE30;
20'b00000110000001001011:ColourData=12'hE30;
20'b00000110010001001011:ColourData=12'hE30;
20'b00000110100001001011:ColourData=12'hF20;
20'b00000110110001001011:ColourData=12'hA70;
20'b00000111000001001011:ColourData=12'h0F0;
20'b00000111010001001011:ColourData=12'h0F0;
20'b00000111100001001011:ColourData=12'h0F0;
20'b00000111110001001011:ColourData=12'h6F6;
20'b00000000000001001100:ColourData=12'h493;
20'b00000000010001001100:ColourData=12'h170;
20'b00000000100001001100:ColourData=12'h170;
20'b00000000110001001100:ColourData=12'h170;
20'b00000001000001001100:ColourData=12'h170;
20'b00000001010001001100:ColourData=12'h170;
20'b00000001100001001100:ColourData=12'h170;
20'b00000001110001001100:ColourData=12'h170;
20'b00000010000001001100:ColourData=12'h170;
20'b00000010010001001100:ColourData=12'h290;
20'b00000010100001001100:ColourData=12'h3D1;
20'b00000010110001001100:ColourData=12'h2A0;
20'b00000011000001001100:ColourData=12'h3D1;
20'b00000011010001001100:ColourData=12'h4F1;
20'b00000011100001001100:ColourData=12'h3D1;
20'b00000011110001001100:ColourData=12'h252;
20'b00000100000001001100:ColourData=12'h0F0;
20'b00000100010001001100:ColourData=12'h3C0;
20'b00000100100001001100:ColourData=12'hB60;
20'b00000100110001001100:ColourData=12'hF20;
20'b00000101000001001100:ColourData=12'hF20;
20'b00000101010001001100:ColourData=12'hF20;
20'b00000101100001001100:ColourData=12'hF20;
20'b00000101110001001100:ColourData=12'hF20;
20'b00000110000001001100:ColourData=12'hF20;
20'b00000110010001001100:ColourData=12'hF20;
20'b00000110100001001100:ColourData=12'hE30;
20'b00000110110001001100:ColourData=12'h790;
20'b00000111000001001100:ColourData=12'h0F0;
20'b00000111010001001100:ColourData=12'h0F0;
20'b00000111100001001100:ColourData=12'h0F0;
20'b00000111110001001100:ColourData=12'h6F6;
20'b00000000000001001101:ColourData=12'h483;
20'b00000000010001001101:ColourData=12'h160;
20'b00000000100001001101:ColourData=12'h160;
20'b00000000110001001101:ColourData=12'h160;
20'b00000001000001001101:ColourData=12'h160;
20'b00000001010001001101:ColourData=12'h160;
20'b00000001100001001101:ColourData=12'h160;
20'b00000001110001001101:ColourData=12'h160;
20'b00000010000001001101:ColourData=12'h170;
20'b00000010010001001101:ColourData=12'h2B1;
20'b00000010100001001101:ColourData=12'h280;
20'b00000010110001001101:ColourData=12'h2B1;
20'b00000011000001001101:ColourData=12'h280;
20'b00000011010001001101:ColourData=12'h3D1;
20'b00000011100001001101:ColourData=12'h2B0;
20'b00000011110001001101:ColourData=12'h252;
20'b00000100000001001101:ColourData=12'h2E0;
20'b00000100010001001101:ColourData=12'hA70;
20'b00000100100001001101:ColourData=12'hA60;
20'b00000100110001001101:ColourData=12'hB50;
20'b00000101000001001101:ColourData=12'hB50;
20'b00000101010001001101:ColourData=12'hC50;
20'b00000101100001001101:ColourData=12'hD40;
20'b00000101110001001101:ColourData=12'hD30;
20'b00000110000001001101:ColourData=12'hE30;
20'b00000110010001001101:ColourData=12'hD40;
20'b00000110100001001101:ColourData=12'h790;
20'b00000110110001001101:ColourData=12'h0F0;
20'b00000111000001001101:ColourData=12'h0F0;
20'b00000111010001001101:ColourData=12'h0F0;
20'b00000111100001001101:ColourData=12'h0F0;
20'b00000111110001001101:ColourData=12'h6F6;
20'b00000000000001001110:ColourData=12'h333;
20'b00000000010001001110:ColourData=12'h000;
20'b00000000100001001110:ColourData=12'h000;
20'b00000000110001001110:ColourData=12'h000;
20'b00000001000001001110:ColourData=12'h000;
20'b00000001010001001110:ColourData=12'h000;
20'b00000001100001001110:ColourData=12'h000;
20'b00000001110001001110:ColourData=12'h000;
20'b00000010000001001110:ColourData=12'h000;
20'b00000010010001001110:ColourData=12'h000;
20'b00000010100001001110:ColourData=12'h000;
20'b00000010110001001110:ColourData=12'h000;
20'b00000011000001001110:ColourData=12'h000;
20'b00000011010001001110:ColourData=12'h000;
20'b00000011100001001110:ColourData=12'h020;
20'b00000011110001001110:ColourData=12'h152;
20'b00000100000001001110:ColourData=12'h1E0;
20'b00000100010001001110:ColourData=12'h790;
20'b00000100100001001110:ColourData=12'h5A0;
20'b00000100110001001110:ColourData=12'h0F0;
20'b00000101000001001110:ColourData=12'h0F0;
20'b00000101010001001110:ColourData=12'h2D0;
20'b00000101100001001110:ColourData=12'hA70;
20'b00000101110001001110:ColourData=12'hA70;
20'b00000110000001001110:ColourData=12'hA70;
20'b00000110010001001110:ColourData=12'h790;
20'b00000110100001001110:ColourData=12'h1E0;
20'b00000110110001001110:ColourData=12'h0F0;
20'b00000111000001001110:ColourData=12'h0F0;
20'b00000111010001001110:ColourData=12'h0F0;
20'b00000111100001001110:ColourData=12'h0F0;
20'b00000111110001001110:ColourData=12'h6F6;
20'b00000000000001001111:ColourData=12'h343;
20'b00000000010001001111:ColourData=12'h000;
20'b00000000100001001111:ColourData=12'h000;
20'b00000000110001001111:ColourData=12'h000;
20'b00000001000001001111:ColourData=12'h000;
20'b00000001010001001111:ColourData=12'h000;
20'b00000001100001001111:ColourData=12'h000;
20'b00000001110001001111:ColourData=12'h000;
20'b00000010000001001111:ColourData=12'h000;
20'b00000010010001001111:ColourData=12'h000;
20'b00000010100001001111:ColourData=12'h000;
20'b00000010110001001111:ColourData=12'h000;
20'b00000011000001001111:ColourData=12'h000;
20'b00000011010001001111:ColourData=12'h020;
20'b00000011100001001111:ColourData=12'h0C0;
20'b00000011110001001111:ColourData=12'h2E2;
20'b00000100000001001111:ColourData=12'h1F0;
20'b00000100010001001111:ColourData=12'h0F0;
20'b00000100100001001111:ColourData=12'h0F0;
20'b00000100110001001111:ColourData=12'h0F0;
20'b00000101000001001111:ColourData=12'h0F0;
20'b00000101010001001111:ColourData=12'h5B0;
20'b00000101100001001111:ColourData=12'hB60;
20'b00000101110001001111:ColourData=12'hB60;
20'b00000110000001001111:ColourData=12'hB60;
20'b00000110010001001111:ColourData=12'hB60;
20'b00000110100001001111:ColourData=12'h790;
20'b00000110110001001111:ColourData=12'h0F0;
20'b00000111000001001111:ColourData=12'h0F0;
20'b00000111010001001111:ColourData=12'h0F0;
20'b00000111100001001111:ColourData=12'h0F0;
20'b00000111110001001111:ColourData=12'h6F6;
20'b00000000000001010000:ColourData=12'h3E3;
20'b00000000010001010000:ColourData=12'h0D0;
20'b00000000100001010000:ColourData=12'h020;
20'b00000000110001010000:ColourData=12'h2A0;
20'b00000001000001010000:ColourData=12'h3E1;
20'b00000001010001010000:ColourData=12'h3D1;
20'b00000001100001010000:ColourData=12'h170;
20'b00000001110001010000:ColourData=12'h170;
20'b00000010000001010000:ColourData=12'h3C1;
20'b00000010010001010000:ColourData=12'h3D1;
20'b00000010100001010000:ColourData=12'h3D1;
20'b00000010110001010000:ColourData=12'h3D1;
20'b00000011000001010000:ColourData=12'h3D1;
20'b00000011010001010000:ColourData=12'h3D1;
20'b00000011100001010000:ColourData=12'h190;
20'b00000011110001010000:ColourData=12'h5F3;
20'b00000100000001010000:ColourData=12'h4F2;
20'b00000100010001010000:ColourData=12'h3F1;
20'b00000100100001010000:ColourData=12'h3F1;
20'b00000100110001010000:ColourData=12'h4E1;
20'b00000101000001010000:ColourData=12'h8A0;
20'b00000101010001010000:ColourData=12'hF30;
20'b00000101100001010000:ColourData=12'hF20;
20'b00000101110001010000:ColourData=12'hE20;
20'b00000110000001010000:ColourData=12'hF20;
20'b00000110010001010000:ColourData=12'hF20;
20'b00000110100001010000:ColourData=12'hC50;
20'b00000110110001010000:ColourData=12'h6C0;
20'b00000111000001010000:ColourData=12'h6C0;
20'b00000111010001010000:ColourData=12'h5D1;
20'b00000111100001010000:ColourData=12'h3F0;
20'b00000111110001010000:ColourData=12'h8F7;
20'b00000000000001010001:ColourData=12'h3F3;
20'b00000000010001010001:ColourData=12'h0F0;
20'b00000000100001010001:ColourData=12'h030;
20'b00000000110001010001:ColourData=12'h3C1;
20'b00000001000001010001:ColourData=12'h4F1;
20'b00000001010001010001:ColourData=12'h3F1;
20'b00000001100001010001:ColourData=12'h280;
20'b00000001110001010001:ColourData=12'h180;
20'b00000010000001010001:ColourData=12'h3E1;
20'b00000010010001010001:ColourData=12'h4F1;
20'b00000010100001010001:ColourData=12'h3F1;
20'b00000010110001010001:ColourData=12'h3F1;
20'b00000011000001010001:ColourData=12'h4F1;
20'b00000011010001010001:ColourData=12'h3E1;
20'b00000011100001010001:ColourData=12'h290;
20'b00000011110001010001:ColourData=12'h5E3;
20'b00000100000001010001:ColourData=12'h4F2;
20'b00000100010001010001:ColourData=12'h3F1;
20'b00000100100001010001:ColourData=12'h3F1;
20'b00000100110001010001:ColourData=12'h6D1;
20'b00000101000001010001:ColourData=12'hD40;
20'b00000101010001010001:ColourData=12'hD30;
20'b00000101100001010001:ColourData=12'hE40;
20'b00000101110001010001:ColourData=12'hF40;
20'b00000110000001010001:ColourData=12'hE40;
20'b00000110010001010001:ColourData=12'hE40;
20'b00000110100001010001:ColourData=12'hF40;
20'b00000110110001010001:ColourData=12'hE50;
20'b00000111000001010001:ColourData=12'hC50;
20'b00000111010001010001:ColourData=12'h990;
20'b00000111100001010001:ColourData=12'h3F1;
20'b00000111110001010001:ColourData=12'h8F7;
20'b00000000000001010010:ColourData=12'h3F3;
20'b00000000010001010010:ColourData=12'h0F0;
20'b00000000100001010010:ColourData=12'h030;
20'b00000000110001010010:ColourData=12'h3C1;
20'b00000001000001010010:ColourData=12'h4F1;
20'b00000001010001010010:ColourData=12'h3F1;
20'b00000001100001010010:ColourData=12'h280;
20'b00000001110001010010:ColourData=12'h170;
20'b00000010000001010010:ColourData=12'h3E1;
20'b00000010010001010010:ColourData=12'h3F1;
20'b00000010100001010010:ColourData=12'h3F1;
20'b00000010110001010010:ColourData=12'h3F1;
20'b00000011000001010010:ColourData=12'h3F1;
20'b00000011010001010010:ColourData=12'h3E1;
20'b00000011100001010010:ColourData=12'h190;
20'b00000011110001010010:ColourData=12'h5E3;
20'b00000100000001010010:ColourData=12'h4F2;
20'b00000100010001010010:ColourData=12'h3F1;
20'b00000100100001010010:ColourData=12'h4F1;
20'b00000100110001010010:ColourData=12'h6C0;
20'b00000101000001010010:ColourData=12'hB70;
20'b00000101010001010010:ColourData=12'hA70;
20'b00000101100001010010:ColourData=12'hC81;
20'b00000101110001010010:ColourData=12'hF93;
20'b00000110000001010010:ColourData=12'hD82;
20'b00000110010001010010:ColourData=12'hB70;
20'b00000110100001010010:ColourData=12'hF93;
20'b00000110110001010010:ColourData=12'hCB2;
20'b00000111000001010010:ColourData=12'h6D1;
20'b00000111010001010010:ColourData=12'h5E1;
20'b00000111100001010010:ColourData=12'h3F0;
20'b00000111110001010010:ColourData=12'h8F7;
20'b00000000000001010011:ColourData=12'h3F3;
20'b00000000010001010011:ColourData=12'h0F0;
20'b00000000100001010011:ColourData=12'h030;
20'b00000000110001010011:ColourData=12'h3C1;
20'b00000001000001010011:ColourData=12'h4F1;
20'b00000001010001010011:ColourData=12'h3F1;
20'b00000001100001010011:ColourData=12'h280;
20'b00000001110001010011:ColourData=12'h170;
20'b00000010000001010011:ColourData=12'h3E1;
20'b00000010010001010011:ColourData=12'h3F1;
20'b00000010100001010011:ColourData=12'h3F1;
20'b00000010110001010011:ColourData=12'h3F1;
20'b00000011000001010011:ColourData=12'h3F1;
20'b00000011010001010011:ColourData=12'h3E1;
20'b00000011100001010011:ColourData=12'h190;
20'b00000011110001010011:ColourData=12'h5E3;
20'b00000100000001010011:ColourData=12'h4F2;
20'b00000100010001010011:ColourData=12'h3F1;
20'b00000100100001010011:ColourData=12'h5D0;
20'b00000100110001010011:ColourData=12'hB80;
20'b00000101000001010011:ColourData=12'hE92;
20'b00000101010001010011:ColourData=12'hB70;
20'b00000101100001010011:ColourData=12'hE92;
20'b00000101110001010011:ColourData=12'hF93;
20'b00000110000001010011:ColourData=12'hE92;
20'b00000110010001010011:ColourData=12'hC81;
20'b00000110100001010011:ColourData=12'hE92;
20'b00000110110001010011:ColourData=12'hF93;
20'b00000111000001010011:ColourData=12'hF93;
20'b00000111010001010011:ColourData=12'hCB3;
20'b00000111100001010011:ColourData=12'h5E1;
20'b00000111110001010011:ColourData=12'h8F7;
20'b00000000000001010100:ColourData=12'h3F3;
20'b00000000010001010100:ColourData=12'h0F0;
20'b00000000100001010100:ColourData=12'h030;
20'b00000000110001010100:ColourData=12'h3C1;
20'b00000001000001010100:ColourData=12'h4F1;
20'b00000001010001010100:ColourData=12'h3F1;
20'b00000001100001010100:ColourData=12'h280;
20'b00000001110001010100:ColourData=12'h170;
20'b00000010000001010100:ColourData=12'h3E1;
20'b00000010010001010100:ColourData=12'h3F1;
20'b00000010100001010100:ColourData=12'h3F1;
20'b00000010110001010100:ColourData=12'h3F1;
20'b00000011000001010100:ColourData=12'h3F1;
20'b00000011010001010100:ColourData=12'h3E1;
20'b00000011100001010100:ColourData=12'h190;
20'b00000011110001010100:ColourData=12'h5E3;
20'b00000100000001010100:ColourData=12'h4F2;
20'b00000100010001010100:ColourData=12'h3F1;
20'b00000100100001010100:ColourData=12'h5D0;
20'b00000100110001010100:ColourData=12'hB70;
20'b00000101000001010100:ColourData=12'hD81;
20'b00000101010001010100:ColourData=12'hB70;
20'b00000101100001010100:ColourData=12'hC81;
20'b00000101110001010100:ColourData=12'hF93;
20'b00000110000001010100:ColourData=12'hF93;
20'b00000110010001010100:ColourData=12'hC81;
20'b00000110100001010100:ColourData=12'hB70;
20'b00000110110001010100:ColourData=12'hE92;
20'b00000111000001010100:ColourData=12'hE82;
20'b00000111010001010100:ColourData=12'hD92;
20'b00000111100001010100:ColourData=12'h8C1;
20'b00000111110001010100:ColourData=12'h8F7;
20'b00000000000001010101:ColourData=12'h3F3;
20'b00000000010001010101:ColourData=12'h0F0;
20'b00000000100001010101:ColourData=12'h030;
20'b00000000110001010101:ColourData=12'h3C1;
20'b00000001000001010101:ColourData=12'h4F1;
20'b00000001010001010101:ColourData=12'h3F1;
20'b00000001100001010101:ColourData=12'h280;
20'b00000001110001010101:ColourData=12'h170;
20'b00000010000001010101:ColourData=12'h3E1;
20'b00000010010001010101:ColourData=12'h3F1;
20'b00000010100001010101:ColourData=12'h3F1;
20'b00000010110001010101:ColourData=12'h3F1;
20'b00000011000001010101:ColourData=12'h3F1;
20'b00000011010001010101:ColourData=12'h3E1;
20'b00000011100001010101:ColourData=12'h190;
20'b00000011110001010101:ColourData=12'h5E3;
20'b00000100000001010101:ColourData=12'h4F2;
20'b00000100010001010101:ColourData=12'h3F1;
20'b00000100100001010101:ColourData=12'h4E1;
20'b00000100110001010101:ColourData=12'h890;
20'b00000101000001010101:ColourData=12'hA90;
20'b00000101010001010101:ColourData=12'hF93;
20'b00000101100001010101:ColourData=12'hF93;
20'b00000101110001010101:ColourData=12'hF93;
20'b00000110000001010101:ColourData=12'hE92;
20'b00000110010001010101:ColourData=12'hB70;
20'b00000110100001010101:ColourData=12'hB70;
20'b00000110110001010101:ColourData=12'hB70;
20'b00000111000001010101:ColourData=12'hA70;
20'b00000111010001010101:ColourData=12'h7B0;
20'b00000111100001010101:ColourData=12'h3F1;
20'b00000111110001010101:ColourData=12'h8F7;
20'b00000000000001010110:ColourData=12'h3F3;
20'b00000000010001010110:ColourData=12'h0F0;
20'b00000000100001010110:ColourData=12'h030;
20'b00000000110001010110:ColourData=12'h3C1;
20'b00000001000001010110:ColourData=12'h4F1;
20'b00000001010001010110:ColourData=12'h3F1;
20'b00000001100001010110:ColourData=12'h280;
20'b00000001110001010110:ColourData=12'h170;
20'b00000010000001010110:ColourData=12'h3E1;
20'b00000010010001010110:ColourData=12'h3F1;
20'b00000010100001010110:ColourData=12'h3F1;
20'b00000010110001010110:ColourData=12'h3F1;
20'b00000011000001010110:ColourData=12'h3F1;
20'b00000011010001010110:ColourData=12'h3E1;
20'b00000011100001010110:ColourData=12'h190;
20'b00000011110001010110:ColourData=12'h5E3;
20'b00000100000001010110:ColourData=12'h4F2;
20'b00000100010001010110:ColourData=12'h3F1;
20'b00000100100001010110:ColourData=12'h3F1;
20'b00000100110001010110:ColourData=12'h3F1;
20'b00000101000001010110:ColourData=12'h7C1;
20'b00000101010001010110:ColourData=12'hE82;
20'b00000101100001010110:ColourData=12'hF82;
20'b00000101110001010110:ColourData=12'hE92;
20'b00000110000001010110:ColourData=12'hE92;
20'b00000110010001010110:ColourData=12'hE92;
20'b00000110100001010110:ColourData=12'hD92;
20'b00000110110001010110:ColourData=12'hCB3;
20'b00000111000001010110:ColourData=12'h9C2;
20'b00000111010001010110:ColourData=12'h3F1;
20'b00000111100001010110:ColourData=12'h3F0;
20'b00000111110001010110:ColourData=12'h8F7;
20'b00000000000001010111:ColourData=12'h3F3;
20'b00000000010001010111:ColourData=12'h0F0;
20'b00000000100001010111:ColourData=12'h030;
20'b00000000110001010111:ColourData=12'h3C1;
20'b00000001000001010111:ColourData=12'h4F1;
20'b00000001010001010111:ColourData=12'h3F1;
20'b00000001100001010111:ColourData=12'h280;
20'b00000001110001010111:ColourData=12'h170;
20'b00000010000001010111:ColourData=12'h3E1;
20'b00000010010001010111:ColourData=12'h3F1;
20'b00000010100001010111:ColourData=12'h3F1;
20'b00000010110001010111:ColourData=12'h3F1;
20'b00000011000001010111:ColourData=12'h3F1;
20'b00000011010001010111:ColourData=12'h3E1;
20'b00000011100001010111:ColourData=12'h190;
20'b00000011110001010111:ColourData=12'h5E3;
20'b00000100000001010111:ColourData=12'h4F2;
20'b00000100010001010111:ColourData=12'h3F1;
20'b00000100100001010111:ColourData=12'h4F1;
20'b00000100110001010111:ColourData=12'h6C0;
20'b00000101000001010111:ColourData=12'hA70;
20'b00000101010001010111:ColourData=12'hB60;
20'b00000101100001010111:ColourData=12'hD40;
20'b00000101110001010111:ColourData=12'hB60;
20'b00000110000001010111:ColourData=12'hB60;
20'b00000110010001010111:ColourData=12'hA70;
20'b00000110100001010111:ColourData=12'h890;
20'b00000110110001010111:ColourData=12'h4E1;
20'b00000111000001010111:ColourData=12'h3F1;
20'b00000111010001010111:ColourData=12'h3F1;
20'b00000111100001010111:ColourData=12'h3F0;
20'b00000111110001010111:ColourData=12'h8F7;
20'b00000000000001011000:ColourData=12'h3F3;
20'b00000000010001011000:ColourData=12'h0F0;
20'b00000000100001011000:ColourData=12'h030;
20'b00000000110001011000:ColourData=12'h3C1;
20'b00000001000001011000:ColourData=12'h4F1;
20'b00000001010001011000:ColourData=12'h3F1;
20'b00000001100001011000:ColourData=12'h280;
20'b00000001110001011000:ColourData=12'h170;
20'b00000010000001011000:ColourData=12'h3E1;
20'b00000010010001011000:ColourData=12'h3F1;
20'b00000010100001011000:ColourData=12'h3F1;
20'b00000010110001011000:ColourData=12'h3F1;
20'b00000011000001011000:ColourData=12'h3F1;
20'b00000011010001011000:ColourData=12'h3E1;
20'b00000011100001011000:ColourData=12'h190;
20'b00000011110001011000:ColourData=12'h5E3;
20'b00000100000001011000:ColourData=12'h4F2;
20'b00000100010001011000:ColourData=12'h3F1;
20'b00000100100001011000:ColourData=12'h5D1;
20'b00000100110001011000:ColourData=12'hA70;
20'b00000101000001011000:ColourData=12'hA70;
20'b00000101010001011000:ColourData=12'hA70;
20'b00000101100001011000:ColourData=12'hC50;
20'b00000101110001011000:ColourData=12'hF30;
20'b00000110000001011000:ColourData=12'hD50;
20'b00000110010001011000:ColourData=12'hB60;
20'b00000110100001011000:ColourData=12'hB60;
20'b00000110110001011000:ColourData=12'h9A1;
20'b00000111000001011000:ColourData=12'h5E1;
20'b00000111010001011000:ColourData=12'h3F1;
20'b00000111100001011000:ColourData=12'h3F0;
20'b00000111110001011000:ColourData=12'h8F7;
20'b00000000000001011001:ColourData=12'h3F3;
20'b00000000010001011001:ColourData=12'h0F0;
20'b00000000100001011001:ColourData=12'h030;
20'b00000000110001011001:ColourData=12'h3C1;
20'b00000001000001011001:ColourData=12'h4F1;
20'b00000001010001011001:ColourData=12'h3F1;
20'b00000001100001011001:ColourData=12'h280;
20'b00000001110001011001:ColourData=12'h170;
20'b00000010000001011001:ColourData=12'h3E1;
20'b00000010010001011001:ColourData=12'h3F1;
20'b00000010100001011001:ColourData=12'h3F1;
20'b00000010110001011001:ColourData=12'h3F1;
20'b00000011000001011001:ColourData=12'h3F1;
20'b00000011010001011001:ColourData=12'h3E1;
20'b00000011100001011001:ColourData=12'h190;
20'b00000011110001011001:ColourData=12'h5E3;
20'b00000100000001011001:ColourData=12'h4F2;
20'b00000100010001011001:ColourData=12'h3F1;
20'b00000100100001011001:ColourData=12'h5D1;
20'b00000100110001011001:ColourData=12'hA70;
20'b00000101000001011001:ColourData=12'hA70;
20'b00000101010001011001:ColourData=12'hB60;
20'b00000101100001011001:ColourData=12'hE30;
20'b00000101110001011001:ColourData=12'hF40;
20'b00000110000001011001:ColourData=12'hF61;
20'b00000110010001011001:ColourData=12'hE20;
20'b00000110100001011001:ColourData=12'hF40;
20'b00000110110001011001:ColourData=12'hF82;
20'b00000111000001011001:ColourData=12'hBA2;
20'b00000111010001011001:ColourData=12'h3F1;
20'b00000111100001011001:ColourData=12'h3F0;
20'b00000111110001011001:ColourData=12'h8F7;
20'b00000000000001011010:ColourData=12'h3F3;
20'b00000000010001011010:ColourData=12'h0F0;
20'b00000000100001011010:ColourData=12'h030;
20'b00000000110001011010:ColourData=12'h3C1;
20'b00000001000001011010:ColourData=12'h4F1;
20'b00000001010001011010:ColourData=12'h3F1;
20'b00000001100001011010:ColourData=12'h280;
20'b00000001110001011010:ColourData=12'h170;
20'b00000010000001011010:ColourData=12'h3E1;
20'b00000010010001011010:ColourData=12'h3F1;
20'b00000010100001011010:ColourData=12'h3F1;
20'b00000010110001011010:ColourData=12'h3F1;
20'b00000011000001011010:ColourData=12'h3F1;
20'b00000011010001011010:ColourData=12'h3E1;
20'b00000011100001011010:ColourData=12'h190;
20'b00000011110001011010:ColourData=12'h5E3;
20'b00000100000001011010:ColourData=12'h4F2;
20'b00000100010001011010:ColourData=12'h3F1;
20'b00000100100001011010:ColourData=12'h5D1;
20'b00000100110001011010:ColourData=12'hB60;
20'b00000101000001011010:ColourData=12'hA70;
20'b00000101010001011010:ColourData=12'hA70;
20'b00000101100001011010:ColourData=12'hC60;
20'b00000101110001011010:ColourData=12'hF40;
20'b00000110000001011010:ColourData=12'hF40;
20'b00000110010001011010:ColourData=12'hF20;
20'b00000110100001011010:ColourData=12'hF30;
20'b00000110110001011010:ColourData=12'hF20;
20'b00000111000001011010:ColourData=12'hB70;
20'b00000111010001011010:ColourData=12'h3F1;
20'b00000111100001011010:ColourData=12'h3F0;
20'b00000111110001011010:ColourData=12'h8F7;
20'b00000000000001011011:ColourData=12'h3F3;
20'b00000000010001011011:ColourData=12'h0F0;
20'b00000000100001011011:ColourData=12'h030;
20'b00000000110001011011:ColourData=12'h3C1;
20'b00000001000001011011:ColourData=12'h4F1;
20'b00000001010001011011:ColourData=12'h3F1;
20'b00000001100001011011:ColourData=12'h280;
20'b00000001110001011011:ColourData=12'h170;
20'b00000010000001011011:ColourData=12'h3E1;
20'b00000010010001011011:ColourData=12'h3F1;
20'b00000010100001011011:ColourData=12'h3F1;
20'b00000010110001011011:ColourData=12'h3F1;
20'b00000011000001011011:ColourData=12'h3F1;
20'b00000011010001011011:ColourData=12'h3E1;
20'b00000011100001011011:ColourData=12'h190;
20'b00000011110001011011:ColourData=12'h5E3;
20'b00000100000001011011:ColourData=12'h4F2;
20'b00000100010001011011:ColourData=12'h3F1;
20'b00000100100001011011:ColourData=12'h5D1;
20'b00000100110001011011:ColourData=12'hC60;
20'b00000101000001011011:ColourData=12'hB60;
20'b00000101010001011011:ColourData=12'hB80;
20'b00000101100001011011:ColourData=12'hFA3;
20'b00000101110001011011:ColourData=12'hF93;
20'b00000110000001011011:ColourData=12'hF61;
20'b00000110010001011011:ColourData=12'hF20;
20'b00000110100001011011:ColourData=12'hF20;
20'b00000110110001011011:ColourData=12'hE30;
20'b00000111000001011011:ColourData=12'h990;
20'b00000111010001011011:ColourData=12'h3F1;
20'b00000111100001011011:ColourData=12'h3F0;
20'b00000111110001011011:ColourData=12'h8F7;
20'b00000000000001011100:ColourData=12'h3F3;
20'b00000000010001011100:ColourData=12'h0F0;
20'b00000000100001011100:ColourData=12'h030;
20'b00000000110001011100:ColourData=12'h3C1;
20'b00000001000001011100:ColourData=12'h4F1;
20'b00000001010001011100:ColourData=12'h3F1;
20'b00000001100001011100:ColourData=12'h280;
20'b00000001110001011100:ColourData=12'h170;
20'b00000010000001011100:ColourData=12'h3E1;
20'b00000010010001011100:ColourData=12'h3F1;
20'b00000010100001011100:ColourData=12'h3F1;
20'b00000010110001011100:ColourData=12'h3F1;
20'b00000011000001011100:ColourData=12'h3F1;
20'b00000011010001011100:ColourData=12'h3E1;
20'b00000011100001011100:ColourData=12'h190;
20'b00000011110001011100:ColourData=12'h5E3;
20'b00000100000001011100:ColourData=12'h4F2;
20'b00000100010001011100:ColourData=12'h3F1;
20'b00000100100001011100:ColourData=12'h3F1;
20'b00000100110001011100:ColourData=12'h5D1;
20'b00000101000001011100:ColourData=12'hB50;
20'b00000101010001011100:ColourData=12'hC60;
20'b00000101100001011100:ColourData=12'hF82;
20'b00000101110001011100:ColourData=12'hF61;
20'b00000110000001011100:ColourData=12'hD40;
20'b00000110010001011100:ColourData=12'hD30;
20'b00000110100001011100:ColourData=12'hE30;
20'b00000110110001011100:ColourData=12'hA70;
20'b00000111000001011100:ColourData=12'h3F1;
20'b00000111010001011100:ColourData=12'h3F1;
20'b00000111100001011100:ColourData=12'h3F0;
20'b00000111110001011100:ColourData=12'h8F7;
20'b00000000000001011101:ColourData=12'h3F3;
20'b00000000010001011101:ColourData=12'h0F0;
20'b00000000100001011101:ColourData=12'h030;
20'b00000000110001011101:ColourData=12'h3C1;
20'b00000001000001011101:ColourData=12'h4F1;
20'b00000001010001011101:ColourData=12'h3F1;
20'b00000001100001011101:ColourData=12'h280;
20'b00000001110001011101:ColourData=12'h170;
20'b00000010000001011101:ColourData=12'h3E1;
20'b00000010010001011101:ColourData=12'h3F1;
20'b00000010100001011101:ColourData=12'h3F1;
20'b00000010110001011101:ColourData=12'h3F1;
20'b00000011000001011101:ColourData=12'h3F1;
20'b00000011010001011101:ColourData=12'h3E1;
20'b00000011100001011101:ColourData=12'h190;
20'b00000011110001011101:ColourData=12'h5E3;
20'b00000100000001011101:ColourData=12'h4F2;
20'b00000100010001011101:ColourData=12'h3F1;
20'b00000100100001011101:ColourData=12'h3F1;
20'b00000100110001011101:ColourData=12'h3F1;
20'b00000101000001011101:ColourData=12'h6C1;
20'b00000101010001011101:ColourData=12'hD40;
20'b00000101100001011101:ColourData=12'hE30;
20'b00000101110001011101:ColourData=12'hC40;
20'b00000110000001011101:ColourData=12'hA70;
20'b00000110010001011101:ColourData=12'hA70;
20'b00000110100001011101:ColourData=12'hA60;
20'b00000110110001011101:ColourData=12'h890;
20'b00000111000001011101:ColourData=12'h4E1;
20'b00000111010001011101:ColourData=12'h3F1;
20'b00000111100001011101:ColourData=12'h3F0;
20'b00000111110001011101:ColourData=12'h8F7;
20'b00000000000001011110:ColourData=12'h3F3;
20'b00000000010001011110:ColourData=12'h0F0;
20'b00000000100001011110:ColourData=12'h030;
20'b00000000110001011110:ColourData=12'h3C1;
20'b00000001000001011110:ColourData=12'h4F1;
20'b00000001010001011110:ColourData=12'h3F1;
20'b00000001100001011110:ColourData=12'h280;
20'b00000001110001011110:ColourData=12'h170;
20'b00000010000001011110:ColourData=12'h3E1;
20'b00000010010001011110:ColourData=12'h3F1;
20'b00000010100001011110:ColourData=12'h3F1;
20'b00000010110001011110:ColourData=12'h3F1;
20'b00000011000001011110:ColourData=12'h3F1;
20'b00000011010001011110:ColourData=12'h3E1;
20'b00000011100001011110:ColourData=12'h290;
20'b00000011110001011110:ColourData=12'h5E3;
20'b00000100000001011110:ColourData=12'h4F2;
20'b00000100010001011110:ColourData=12'h3F1;
20'b00000100100001011110:ColourData=12'h3F1;
20'b00000100110001011110:ColourData=12'h3F1;
20'b00000101000001011110:ColourData=12'h5D1;
20'b00000101010001011110:ColourData=12'hA70;
20'b00000101100001011110:ColourData=12'hA70;
20'b00000101110001011110:ColourData=12'hA70;
20'b00000110000001011110:ColourData=12'hA70;
20'b00000110010001011110:ColourData=12'h980;
20'b00000110100001011110:ColourData=12'h890;
20'b00000110110001011110:ColourData=12'h880;
20'b00000111000001011110:ColourData=12'h7B0;
20'b00000111010001011110:ColourData=12'h3F1;
20'b00000111100001011110:ColourData=12'h3F0;
20'b00000111110001011110:ColourData=12'h8F7;
20'b00000000000001011111:ColourData=12'h3E3;
20'b00000000010001011111:ColourData=12'h0E0;
20'b00000000100001011111:ColourData=12'h030;
20'b00000000110001011111:ColourData=12'h2B1;
20'b00000001000001011111:ColourData=12'h3E1;
20'b00000001010001011111:ColourData=12'h3E1;
20'b00000001100001011111:ColourData=12'h180;
20'b00000001110001011111:ColourData=12'h170;
20'b00000010000001011111:ColourData=12'h3E1;
20'b00000010010001011111:ColourData=12'h3E1;
20'b00000010100001011111:ColourData=12'h3F1;
20'b00000010110001011111:ColourData=12'h3F1;
20'b00000011000001011111:ColourData=12'h3F1;
20'b00000011010001011111:ColourData=12'h3D1;
20'b00000011100001011111:ColourData=12'h190;
20'b00000011110001011111:ColourData=12'h5E3;
20'b00000100000001011111:ColourData=12'h4F2;
20'b00000100010001011111:ColourData=12'h3F1;
20'b00000100100001011111:ColourData=12'h3F1;
20'b00000100110001011111:ColourData=12'h3F1;
20'b00000101000001011111:ColourData=12'h5D1;
20'b00000101010001011111:ColourData=12'hB60;
20'b00000101100001011111:ColourData=12'hB60;
20'b00000101110001011111:ColourData=12'hB60;
20'b00000110000001011111:ColourData=12'hB60;
20'b00000110010001011111:ColourData=12'h980;
20'b00000110100001011111:ColourData=12'h5D1;
20'b00000110110001011111:ColourData=12'h3F1;
20'b00000111000001011111:ColourData=12'h3F1;
20'b00000111010001011111:ColourData=12'h3F1;
20'b00000111100001011111:ColourData=12'h3F0;
20'b00000111110001011111:ColourData=12'h8F7;
20'b00000000000001100000:ColourData=12'h493;
20'b00000000010001100000:ColourData=12'h180;
20'b00000000100001100000:ColourData=12'h170;
20'b00000000110001100000:ColourData=12'h180;
20'b00000001000001100000:ColourData=12'h180;
20'b00000001010001100000:ColourData=12'h180;
20'b00000001100001100000:ColourData=12'h170;
20'b00000001110001100000:ColourData=12'h180;
20'b00000010000001100000:ColourData=12'h3D1;
20'b00000010010001100000:ColourData=12'h2A0;
20'b00000010100001100000:ColourData=12'h3D1;
20'b00000010110001100000:ColourData=12'h3F1;
20'b00000011000001100000:ColourData=12'h3D1;
20'b00000011010001100000:ColourData=12'h030;
20'b00000011100001100000:ColourData=12'h0D0;
20'b00000011110001100000:ColourData=12'h2F2;
20'b00000100000001100000:ColourData=12'h4F2;
20'b00000100010001100000:ColourData=12'h3F1;
20'b00000100100001100000:ColourData=12'h3F1;
20'b00000100110001100000:ColourData=12'h4E1;
20'b00000101000001100000:ColourData=12'h8A0;
20'b00000101010001100000:ColourData=12'hF20;
20'b00000101100001100000:ColourData=12'hF20;
20'b00000101110001100000:ColourData=12'hE20;
20'b00000110000001100000:ColourData=12'hF20;
20'b00000110010001100000:ColourData=12'hF20;
20'b00000110100001100000:ColourData=12'hC60;
20'b00000110110001100000:ColourData=12'h6C1;
20'b00000111000001100000:ColourData=12'h6C1;
20'b00000111010001100000:ColourData=12'h5D1;
20'b00000111100001100000:ColourData=12'h3F0;
20'b00000111110001100000:ColourData=12'h8F7;
20'b00000000000001100001:ColourData=12'h493;
20'b00000000010001100001:ColourData=12'h170;
20'b00000000100001100001:ColourData=12'h170;
20'b00000000110001100001:ColourData=12'h170;
20'b00000001000001100001:ColourData=12'h170;
20'b00000001010001100001:ColourData=12'h170;
20'b00000001100001100001:ColourData=12'h170;
20'b00000001110001100001:ColourData=12'h170;
20'b00000010000001100001:ColourData=12'h290;
20'b00000010010001100001:ColourData=12'h3C1;
20'b00000010100001100001:ColourData=12'h2A0;
20'b00000010110001100001:ColourData=12'h3E1;
20'b00000011000001100001:ColourData=12'h3D1;
20'b00000011010001100001:ColourData=12'h020;
20'b00000011100001100001:ColourData=12'h0E0;
20'b00000011110001100001:ColourData=12'h2F2;
20'b00000100000001100001:ColourData=12'h4F2;
20'b00000100010001100001:ColourData=12'h3F1;
20'b00000100100001100001:ColourData=12'h3F1;
20'b00000100110001100001:ColourData=12'h6D1;
20'b00000101000001100001:ColourData=12'hD40;
20'b00000101010001100001:ColourData=12'hD30;
20'b00000101100001100001:ColourData=12'hE40;
20'b00000101110001100001:ColourData=12'hF40;
20'b00000110000001100001:ColourData=12'hE40;
20'b00000110010001100001:ColourData=12'hE40;
20'b00000110100001100001:ColourData=12'hF40;
20'b00000110110001100001:ColourData=12'hE50;
20'b00000111000001100001:ColourData=12'hC50;
20'b00000111010001100001:ColourData=12'h990;
20'b00000111100001100001:ColourData=12'h3F1;
20'b00000111110001100001:ColourData=12'h8F7;
20'b00000000000001100010:ColourData=12'h493;
20'b00000000010001100010:ColourData=12'h170;
20'b00000000100001100010:ColourData=12'h170;
20'b00000000110001100010:ColourData=12'h170;
20'b00000001000001100010:ColourData=12'h170;
20'b00000001010001100010:ColourData=12'h170;
20'b00000001100001100010:ColourData=12'h170;
20'b00000001110001100010:ColourData=12'h180;
20'b00000010000001100010:ColourData=12'h3C1;
20'b00000010010001100010:ColourData=12'h2A0;
20'b00000010100001100010:ColourData=12'h3D1;
20'b00000010110001100010:ColourData=12'h3F1;
20'b00000011000001100010:ColourData=12'h3D1;
20'b00000011010001100010:ColourData=12'h020;
20'b00000011100001100010:ColourData=12'h0D0;
20'b00000011110001100010:ColourData=12'h2F2;
20'b00000100000001100010:ColourData=12'h4F2;
20'b00000100010001100010:ColourData=12'h3F1;
20'b00000100100001100010:ColourData=12'h4F1;
20'b00000100110001100010:ColourData=12'h6C0;
20'b00000101000001100010:ColourData=12'hB70;
20'b00000101010001100010:ColourData=12'hA70;
20'b00000101100001100010:ColourData=12'hC81;
20'b00000101110001100010:ColourData=12'hF93;
20'b00000110000001100010:ColourData=12'hD82;
20'b00000110010001100010:ColourData=12'hB70;
20'b00000110100001100010:ColourData=12'hF93;
20'b00000110110001100010:ColourData=12'hCB2;
20'b00000111000001100010:ColourData=12'h6D1;
20'b00000111010001100010:ColourData=12'h5E1;
20'b00000111100001100010:ColourData=12'h3F0;
20'b00000111110001100010:ColourData=12'h8F7;
20'b00000000000001100011:ColourData=12'h493;
20'b00000000010001100011:ColourData=12'h170;
20'b00000000100001100011:ColourData=12'h170;
20'b00000000110001100011:ColourData=12'h170;
20'b00000001000001100011:ColourData=12'h170;
20'b00000001010001100011:ColourData=12'h170;
20'b00000001100001100011:ColourData=12'h170;
20'b00000001110001100011:ColourData=12'h170;
20'b00000010000001100011:ColourData=12'h290;
20'b00000010010001100011:ColourData=12'h3C1;
20'b00000010100001100011:ColourData=12'h2A0;
20'b00000010110001100011:ColourData=12'h3E1;
20'b00000011000001100011:ColourData=12'h3D1;
20'b00000011010001100011:ColourData=12'h020;
20'b00000011100001100011:ColourData=12'h0D0;
20'b00000011110001100011:ColourData=12'h2F2;
20'b00000100000001100011:ColourData=12'h4F2;
20'b00000100010001100011:ColourData=12'h3F1;
20'b00000100100001100011:ColourData=12'h5D0;
20'b00000100110001100011:ColourData=12'hB80;
20'b00000101000001100011:ColourData=12'hE92;
20'b00000101010001100011:ColourData=12'hB70;
20'b00000101100001100011:ColourData=12'hE92;
20'b00000101110001100011:ColourData=12'hF93;
20'b00000110000001100011:ColourData=12'hE92;
20'b00000110010001100011:ColourData=12'hC81;
20'b00000110100001100011:ColourData=12'hE92;
20'b00000110110001100011:ColourData=12'hF93;
20'b00000111000001100011:ColourData=12'hF93;
20'b00000111010001100011:ColourData=12'hCB3;
20'b00000111100001100011:ColourData=12'h5E1;
20'b00000111110001100011:ColourData=12'h8F7;
20'b00000000000001100100:ColourData=12'h493;
20'b00000000010001100100:ColourData=12'h170;
20'b00000000100001100100:ColourData=12'h170;
20'b00000000110001100100:ColourData=12'h170;
20'b00000001000001100100:ColourData=12'h170;
20'b00000001010001100100:ColourData=12'h170;
20'b00000001100001100100:ColourData=12'h170;
20'b00000001110001100100:ColourData=12'h180;
20'b00000010000001100100:ColourData=12'h3C1;
20'b00000010010001100100:ColourData=12'h2A0;
20'b00000010100001100100:ColourData=12'h3D1;
20'b00000010110001100100:ColourData=12'h3F1;
20'b00000011000001100100:ColourData=12'h3D1;
20'b00000011010001100100:ColourData=12'h020;
20'b00000011100001100100:ColourData=12'h0D0;
20'b00000011110001100100:ColourData=12'h2F2;
20'b00000100000001100100:ColourData=12'h4F2;
20'b00000100010001100100:ColourData=12'h3F1;
20'b00000100100001100100:ColourData=12'h5D0;
20'b00000100110001100100:ColourData=12'hB70;
20'b00000101000001100100:ColourData=12'hD81;
20'b00000101010001100100:ColourData=12'hB70;
20'b00000101100001100100:ColourData=12'hC81;
20'b00000101110001100100:ColourData=12'hF93;
20'b00000110000001100100:ColourData=12'hF93;
20'b00000110010001100100:ColourData=12'hC81;
20'b00000110100001100100:ColourData=12'hB70;
20'b00000110110001100100:ColourData=12'hE92;
20'b00000111000001100100:ColourData=12'hE82;
20'b00000111010001100100:ColourData=12'hD92;
20'b00000111100001100100:ColourData=12'h8C1;
20'b00000111110001100100:ColourData=12'h8F7;
20'b00000000000001100101:ColourData=12'h493;
20'b00000000010001100101:ColourData=12'h170;
20'b00000000100001100101:ColourData=12'h170;
20'b00000000110001100101:ColourData=12'h170;
20'b00000001000001100101:ColourData=12'h170;
20'b00000001010001100101:ColourData=12'h170;
20'b00000001100001100101:ColourData=12'h170;
20'b00000001110001100101:ColourData=12'h170;
20'b00000010000001100101:ColourData=12'h290;
20'b00000010010001100101:ColourData=12'h3C1;
20'b00000010100001100101:ColourData=12'h2A0;
20'b00000010110001100101:ColourData=12'h3E1;
20'b00000011000001100101:ColourData=12'h3D1;
20'b00000011010001100101:ColourData=12'h020;
20'b00000011100001100101:ColourData=12'h0D0;
20'b00000011110001100101:ColourData=12'h2F2;
20'b00000100000001100101:ColourData=12'h4F2;
20'b00000100010001100101:ColourData=12'h3F1;
20'b00000100100001100101:ColourData=12'h4E1;
20'b00000100110001100101:ColourData=12'h890;
20'b00000101000001100101:ColourData=12'hA90;
20'b00000101010001100101:ColourData=12'hF93;
20'b00000101100001100101:ColourData=12'hF93;
20'b00000101110001100101:ColourData=12'hF93;
20'b00000110000001100101:ColourData=12'hE92;
20'b00000110010001100101:ColourData=12'hB70;
20'b00000110100001100101:ColourData=12'hB70;
20'b00000110110001100101:ColourData=12'hB70;
20'b00000111000001100101:ColourData=12'hA70;
20'b00000111010001100101:ColourData=12'h7B0;
20'b00000111100001100101:ColourData=12'h3F1;
20'b00000111110001100101:ColourData=12'h8F7;
20'b00000000000001100110:ColourData=12'h493;
20'b00000000010001100110:ColourData=12'h170;
20'b00000000100001100110:ColourData=12'h170;
20'b00000000110001100110:ColourData=12'h170;
20'b00000001000001100110:ColourData=12'h170;
20'b00000001010001100110:ColourData=12'h170;
20'b00000001100001100110:ColourData=12'h170;
20'b00000001110001100110:ColourData=12'h180;
20'b00000010000001100110:ColourData=12'h3C1;
20'b00000010010001100110:ColourData=12'h2A0;
20'b00000010100001100110:ColourData=12'h3D1;
20'b00000010110001100110:ColourData=12'h3F1;
20'b00000011000001100110:ColourData=12'h3D1;
20'b00000011010001100110:ColourData=12'h020;
20'b00000011100001100110:ColourData=12'h0D0;
20'b00000011110001100110:ColourData=12'h2F2;
20'b00000100000001100110:ColourData=12'h4F2;
20'b00000100010001100110:ColourData=12'h3F1;
20'b00000100100001100110:ColourData=12'h5D1;
20'b00000100110001100110:ColourData=12'h5D0;
20'b00000101000001100110:ColourData=12'h7C1;
20'b00000101010001100110:ColourData=12'hE82;
20'b00000101100001100110:ColourData=12'hF82;
20'b00000101110001100110:ColourData=12'hF82;
20'b00000110000001100110:ColourData=12'hE92;
20'b00000110010001100110:ColourData=12'hE92;
20'b00000110100001100110:ColourData=12'hD92;
20'b00000110110001100110:ColourData=12'hCB3;
20'b00000111000001100110:ColourData=12'h9C2;
20'b00000111010001100110:ColourData=12'h3F1;
20'b00000111100001100110:ColourData=12'h3F0;
20'b00000111110001100110:ColourData=12'h8F7;
20'b00000000000001100111:ColourData=12'h493;
20'b00000000010001100111:ColourData=12'h170;
20'b00000000100001100111:ColourData=12'h170;
20'b00000000110001100111:ColourData=12'h170;
20'b00000001000001100111:ColourData=12'h170;
20'b00000001010001100111:ColourData=12'h170;
20'b00000001100001100111:ColourData=12'h170;
20'b00000001110001100111:ColourData=12'h170;
20'b00000010000001100111:ColourData=12'h290;
20'b00000010010001100111:ColourData=12'h3C1;
20'b00000010100001100111:ColourData=12'h2A0;
20'b00000010110001100111:ColourData=12'h3E1;
20'b00000011000001100111:ColourData=12'h3D1;
20'b00000011010001100111:ColourData=12'h020;
20'b00000011100001100111:ColourData=12'h0D0;
20'b00000011110001100111:ColourData=12'h2F2;
20'b00000100000001100111:ColourData=12'h6E2;
20'b00000100010001100111:ColourData=12'h7C1;
20'b00000100100001100111:ColourData=12'h970;
20'b00000100110001100111:ColourData=12'hA70;
20'b00000101000001100111:ColourData=12'hA70;
20'b00000101010001100111:ColourData=12'hB60;
20'b00000101100001100111:ColourData=12'hF20;
20'b00000101110001100111:ColourData=12'hE30;
20'b00000110000001100111:ColourData=12'hB60;
20'b00000110010001100111:ColourData=12'hA70;
20'b00000110100001100111:ColourData=12'h890;
20'b00000110110001100111:ColourData=12'h5D1;
20'b00000111000001100111:ColourData=12'h6E2;
20'b00000111010001100111:ColourData=12'h6E1;
20'b00000111100001100111:ColourData=12'h6E1;
20'b00000111110001100111:ColourData=12'hAE7;
20'b00000000000001101000:ColourData=12'h493;
20'b00000000010001101000:ColourData=12'h170;
20'b00000000100001101000:ColourData=12'h170;
20'b00000000110001101000:ColourData=12'h170;
20'b00000001000001101000:ColourData=12'h170;
20'b00000001010001101000:ColourData=12'h170;
20'b00000001100001101000:ColourData=12'h170;
20'b00000001110001101000:ColourData=12'h180;
20'b00000010000001101000:ColourData=12'h3C1;
20'b00000010010001101000:ColourData=12'h2A0;
20'b00000010100001101000:ColourData=12'h3D1;
20'b00000010110001101000:ColourData=12'h3F1;
20'b00000011000001101000:ColourData=12'h3D1;
20'b00000011010001101000:ColourData=12'h020;
20'b00000011100001101000:ColourData=12'h0E0;
20'b00000011110001101000:ColourData=12'h3E2;
20'b00000100000001101000:ColourData=12'hFA4;
20'b00000100010001101000:ColourData=12'hE92;
20'b00000100100001101000:ColourData=12'hB70;
20'b00000100110001101000:ColourData=12'hB70;
20'b00000101000001101000:ColourData=12'hA70;
20'b00000101010001101000:ColourData=12'hB60;
20'b00000101100001101000:ColourData=12'hF30;
20'b00000101110001101000:ColourData=12'hF40;
20'b00000110000001101000:ColourData=12'hD30;
20'b00000110010001101000:ColourData=12'hB60;
20'b00000110100001101000:ColourData=12'hA60;
20'b00000110110001101000:ColourData=12'hB80;
20'b00000111000001101000:ColourData=12'hE92;
20'b00000111010001101000:ColourData=12'hF93;
20'b00000111100001101000:ColourData=12'hF93;
20'b00000111110001101000:ColourData=12'hFC8;
20'b00000000000001101001:ColourData=12'h493;
20'b00000000010001101001:ColourData=12'h170;
20'b00000000100001101001:ColourData=12'h170;
20'b00000000110001101001:ColourData=12'h170;
20'b00000001000001101001:ColourData=12'h170;
20'b00000001010001101001:ColourData=12'h170;
20'b00000001100001101001:ColourData=12'h170;
20'b00000001110001101001:ColourData=12'h170;
20'b00000010000001101001:ColourData=12'h290;
20'b00000010010001101001:ColourData=12'h3C1;
20'b00000010100001101001:ColourData=12'h2A0;
20'b00000010110001101001:ColourData=12'h3E1;
20'b00000011000001101001:ColourData=12'h3D1;
20'b00000011010001101001:ColourData=12'h020;
20'b00000011100001101001:ColourData=12'h0E0;
20'b00000011110001101001:ColourData=12'h4E2;
20'b00000100000001101001:ColourData=12'hF94;
20'b00000100010001101001:ColourData=12'hF93;
20'b00000100100001101001:ColourData=12'hEA3;
20'b00000100110001101001:ColourData=12'hCA2;
20'b00000101000001101001:ColourData=12'hB60;
20'b00000101010001101001:ColourData=12'hC50;
20'b00000101100001101001:ColourData=12'hF40;
20'b00000101110001101001:ColourData=12'hF61;
20'b00000110000001101001:ColourData=12'hF20;
20'b00000110010001101001:ColourData=12'hF20;
20'b00000110100001101001:ColourData=12'hD30;
20'b00000110110001101001:ColourData=12'hA70;
20'b00000111000001101001:ColourData=12'hA90;
20'b00000111010001101001:ColourData=12'hE92;
20'b00000111100001101001:ColourData=12'hD92;
20'b00000111110001101001:ColourData=12'hDC8;
20'b00000000000001101010:ColourData=12'h493;
20'b00000000010001101010:ColourData=12'h170;
20'b00000000100001101010:ColourData=12'h170;
20'b00000000110001101010:ColourData=12'h170;
20'b00000001000001101010:ColourData=12'h170;
20'b00000001010001101010:ColourData=12'h170;
20'b00000001100001101010:ColourData=12'h170;
20'b00000001110001101010:ColourData=12'h180;
20'b00000010000001101010:ColourData=12'h3C1;
20'b00000010010001101010:ColourData=12'h2A0;
20'b00000010100001101010:ColourData=12'h3D1;
20'b00000010110001101010:ColourData=12'h3F1;
20'b00000011000001101010:ColourData=12'h3D1;
20'b00000011010001101010:ColourData=12'h020;
20'b00000011100001101010:ColourData=12'h0E0;
20'b00000011110001101010:ColourData=12'h3F2;
20'b00000100000001101010:ColourData=12'hCB3;
20'b00000100010001101010:ColourData=12'hCB3;
20'b00000100100001101010:ColourData=12'hBB2;
20'b00000100110001101010:ColourData=12'h8A0;
20'b00000101000001101010:ColourData=12'hE30;
20'b00000101010001101010:ColourData=12'hF30;
20'b00000101100001101010:ColourData=12'hF30;
20'b00000101110001101010:ColourData=12'hF30;
20'b00000110000001101010:ColourData=12'hF30;
20'b00000110010001101010:ColourData=12'hF30;
20'b00000110100001101010:ColourData=12'hF20;
20'b00000110110001101010:ColourData=12'hB60;
20'b00000111000001101010:ColourData=12'h6B0;
20'b00000111010001101010:ColourData=12'hA60;
20'b00000111100001101010:ColourData=12'h7A0;
20'b00000111110001101010:ColourData=12'h8F7;
20'b00000000000001101011:ColourData=12'h493;
20'b00000000010001101011:ColourData=12'h170;
20'b00000000100001101011:ColourData=12'h170;
20'b00000000110001101011:ColourData=12'h170;
20'b00000001000001101011:ColourData=12'h170;
20'b00000001010001101011:ColourData=12'h170;
20'b00000001100001101011:ColourData=12'h170;
20'b00000001110001101011:ColourData=12'h170;
20'b00000010000001101011:ColourData=12'h290;
20'b00000010010001101011:ColourData=12'h3C1;
20'b00000010100001101011:ColourData=12'h2A0;
20'b00000010110001101011:ColourData=12'h3E1;
20'b00000011000001101011:ColourData=12'h3D1;
20'b00000011010001101011:ColourData=12'h020;
20'b00000011100001101011:ColourData=12'h0D0;
20'b00000011110001101011:ColourData=12'h2F2;
20'b00000100000001101011:ColourData=12'h4F2;
20'b00000100010001101011:ColourData=12'h4F1;
20'b00000100100001101011:ColourData=12'h8A0;
20'b00000100110001101011:ColourData=12'hE30;
20'b00000101000001101011:ColourData=12'hF20;
20'b00000101010001101011:ColourData=12'hF30;
20'b00000101100001101011:ColourData=12'hF20;
20'b00000101110001101011:ColourData=12'hF20;
20'b00000110000001101011:ColourData=12'hF20;
20'b00000110010001101011:ColourData=12'hF30;
20'b00000110100001101011:ColourData=12'hF20;
20'b00000110110001101011:ColourData=12'hD40;
20'b00000111000001101011:ColourData=12'hA70;
20'b00000111010001101011:ColourData=12'hA60;
20'b00000111100001101011:ColourData=12'h7A0;
20'b00000111110001101011:ColourData=12'h8F7;
20'b00000000000001101100:ColourData=12'h493;
20'b00000000010001101100:ColourData=12'h170;
20'b00000000100001101100:ColourData=12'h170;
20'b00000000110001101100:ColourData=12'h170;
20'b00000001000001101100:ColourData=12'h170;
20'b00000001010001101100:ColourData=12'h170;
20'b00000001100001101100:ColourData=12'h170;
20'b00000001110001101100:ColourData=12'h180;
20'b00000010000001101100:ColourData=12'h3C1;
20'b00000010010001101100:ColourData=12'h2A0;
20'b00000010100001101100:ColourData=12'h3D1;
20'b00000010110001101100:ColourData=12'h3F1;
20'b00000011000001101100:ColourData=12'h3D1;
20'b00000011010001101100:ColourData=12'h020;
20'b00000011100001101100:ColourData=12'h0D0;
20'b00000011110001101100:ColourData=12'h2F2;
20'b00000100000001101100:ColourData=12'h4F2;
20'b00000100010001101100:ColourData=12'h6B0;
20'b00000100100001101100:ColourData=12'hD30;
20'b00000100110001101100:ColourData=12'hF20;
20'b00000101000001101100:ColourData=12'hF20;
20'b00000101010001101100:ColourData=12'hF20;
20'b00000101100001101100:ColourData=12'hE30;
20'b00000101110001101100:ColourData=12'hC50;
20'b00000110000001101100:ColourData=12'hD40;
20'b00000110010001101100:ColourData=12'hF20;
20'b00000110100001101100:ColourData=12'hF20;
20'b00000110110001101100:ColourData=12'hD40;
20'b00000111000001101100:ColourData=12'hA70;
20'b00000111010001101100:ColourData=12'hA60;
20'b00000111100001101100:ColourData=12'h7A0;
20'b00000111110001101100:ColourData=12'h8F7;
20'b00000000000001101101:ColourData=12'h493;
20'b00000000010001101101:ColourData=12'h170;
20'b00000000100001101101:ColourData=12'h170;
20'b00000000110001101101:ColourData=12'h170;
20'b00000001000001101101:ColourData=12'h170;
20'b00000001010001101101:ColourData=12'h170;
20'b00000001100001101101:ColourData=12'h170;
20'b00000001110001101101:ColourData=12'h170;
20'b00000010000001101101:ColourData=12'h290;
20'b00000010010001101101:ColourData=12'h3C1;
20'b00000010100001101101:ColourData=12'h2A0;
20'b00000010110001101101:ColourData=12'h3E1;
20'b00000011000001101101:ColourData=12'h3D1;
20'b00000011010001101101:ColourData=12'h020;
20'b00000011100001101101:ColourData=12'h0D0;
20'b00000011110001101101:ColourData=12'h2F2;
20'b00000100000001101101:ColourData=12'h5D1;
20'b00000100010001101101:ColourData=12'hA70;
20'b00000100100001101101:ColourData=12'hB60;
20'b00000100110001101101:ColourData=12'hD30;
20'b00000101000001101101:ColourData=12'hD40;
20'b00000101010001101101:ColourData=12'hC50;
20'b00000101100001101101:ColourData=12'hA80;
20'b00000101110001101101:ColourData=12'h3F1;
20'b00000110000001101101:ColourData=12'h6C1;
20'b00000110010001101101:ColourData=12'hC50;
20'b00000110100001101101:ColourData=12'hC50;
20'b00000110110001101101:ColourData=12'hB60;
20'b00000111000001101101:ColourData=12'h890;
20'b00000111010001101101:ColourData=12'h880;
20'b00000111100001101101:ColourData=12'h6B0;
20'b00000111110001101101:ColourData=12'h8F7;
20'b00000000000001101110:ColourData=12'h493;
20'b00000000010001101110:ColourData=12'h170;
20'b00000000100001101110:ColourData=12'h170;
20'b00000000110001101110:ColourData=12'h170;
20'b00000001000001101110:ColourData=12'h170;
20'b00000001010001101110:ColourData=12'h170;
20'b00000001100001101110:ColourData=12'h170;
20'b00000001110001101110:ColourData=12'h170;
20'b00000010000001101110:ColourData=12'h3C1;
20'b00000010010001101110:ColourData=12'h2A0;
20'b00000010100001101110:ColourData=12'h3D1;
20'b00000010110001101110:ColourData=12'h4F1;
20'b00000011000001101110:ColourData=12'h3D1;
20'b00000011010001101110:ColourData=12'h020;
20'b00000011100001101110:ColourData=12'h0D0;
20'b00000011110001101110:ColourData=12'h2F2;
20'b00000100000001101110:ColourData=12'h5E2;
20'b00000100010001101110:ColourData=12'h880;
20'b00000100100001101110:ColourData=12'hA70;
20'b00000100110001101110:ColourData=12'hA60;
20'b00000101000001101110:ColourData=12'h980;
20'b00000101010001101110:ColourData=12'h5D1;
20'b00000101100001101110:ColourData=12'h3F1;
20'b00000101110001101110:ColourData=12'h3F1;
20'b00000110000001101110:ColourData=12'h3F1;
20'b00000110010001101110:ColourData=12'h3F1;
20'b00000110100001101110:ColourData=12'h3F1;
20'b00000110110001101110:ColourData=12'h3F1;
20'b00000111000001101110:ColourData=12'h3F1;
20'b00000111010001101110:ColourData=12'h3F1;
20'b00000111100001101110:ColourData=12'h3F0;
20'b00000111110001101110:ColourData=12'h8F7;
20'b00000000000001101111:ColourData=12'h493;
20'b00000000010001101111:ColourData=12'h180;
20'b00000000100001101111:ColourData=12'h180;
20'b00000000110001101111:ColourData=12'h180;
20'b00000001000001101111:ColourData=12'h180;
20'b00000001010001101111:ColourData=12'h180;
20'b00000001100001101111:ColourData=12'h180;
20'b00000001110001101111:ColourData=12'h180;
20'b00000010000001101111:ColourData=12'h290;
20'b00000010010001101111:ColourData=12'h2D1;
20'b00000010100001101111:ColourData=12'h2A0;
20'b00000010110001101111:ColourData=12'h3E1;
20'b00000011000001101111:ColourData=12'h3D1;
20'b00000011010001101111:ColourData=12'h030;
20'b00000011100001101111:ColourData=12'h0E0;
20'b00000011110001101111:ColourData=12'h2F2;
20'b00000100000001101111:ColourData=12'h4F2;
20'b00000100010001101111:ColourData=12'h4E1;
20'b00000100100001101111:ColourData=12'h890;
20'b00000100110001101111:ColourData=12'h890;
20'b00000101000001101111:ColourData=12'h890;
20'b00000101010001101111:ColourData=12'h7A0;
20'b00000101100001101111:ColourData=12'h6C1;
20'b00000101110001101111:ColourData=12'h6C1;
20'b00000110000001101111:ColourData=12'h6C1;
20'b00000110010001101111:ColourData=12'h6C1;
20'b00000110100001101111:ColourData=12'h6C1;
20'b00000110110001101111:ColourData=12'h5D1;
20'b00000111000001101111:ColourData=12'h3F1;
20'b00000111010001101111:ColourData=12'h3F1;
20'b00000111100001101111:ColourData=12'h3F0;
20'b00000111110001101111:ColourData=12'h8F7;
20'b00000000000001110000:ColourData=12'h3E3;
20'b00000000010001110000:ColourData=12'h0E0;
20'b00000000100001110000:ColourData=12'h0E0;
20'b00000000110001110000:ColourData=12'h0E0;
20'b00000001000001110000:ColourData=12'h0E0;
20'b00000001010001110000:ColourData=12'h0E0;
20'b00000001100001110000:ColourData=12'h0E0;
20'b00000001110001110000:ColourData=12'h3E1;
20'b00000010000001110000:ColourData=12'h3E1;
20'b00000010010001110000:ColourData=12'h0F0;
20'b00000010100001110000:ColourData=12'h0E0;
20'b00000010110001110000:ColourData=12'h0F0;
20'b00000011000001110000:ColourData=12'h0F0;
20'b00000011010001110000:ColourData=12'h0E0;
20'b00000011100001110000:ColourData=12'h0F0;
20'b00000011110001110000:ColourData=12'h2F2;
20'b00000100000001110000:ColourData=12'h4F2;
20'b00000100010001110000:ColourData=12'h3F1;
20'b00000100100001110000:ColourData=12'h3F1;
20'b00000100110001110000:ColourData=12'h4F1;
20'b00000101000001110000:ColourData=12'h5D1;
20'b00000101010001110000:ColourData=12'h890;
20'b00000101100001110000:ColourData=12'hF30;
20'b00000101110001110000:ColourData=12'hF20;
20'b00000110000001110000:ColourData=12'hF30;
20'b00000110010001110000:ColourData=12'hE20;
20'b00000110100001110000:ColourData=12'hF20;
20'b00000110110001110000:ColourData=12'hC60;
20'b00000111000001110000:ColourData=12'h6C0;
20'b00000111010001110000:ColourData=12'h5D1;
20'b00000111100001110000:ColourData=12'h3F0;
20'b00000111110001110000:ColourData=12'h8F7;
20'b00000000000001110001:ColourData=12'h3F3;
20'b00000000010001110001:ColourData=12'h0F0;
20'b00000000100001110001:ColourData=12'h0F0;
20'b00000000110001110001:ColourData=12'h0F0;
20'b00000001000001110001:ColourData=12'h0F0;
20'b00000001010001110001:ColourData=12'h0F0;
20'b00000001100001110001:ColourData=12'h0F0;
20'b00000001110001110001:ColourData=12'h3F1;
20'b00000010000001110001:ColourData=12'h3F1;
20'b00000010010001110001:ColourData=12'h0F0;
20'b00000010100001110001:ColourData=12'h0F0;
20'b00000010110001110001:ColourData=12'h0F0;
20'b00000011000001110001:ColourData=12'h0F0;
20'b00000011010001110001:ColourData=12'h0F0;
20'b00000011100001110001:ColourData=12'h0F0;
20'b00000011110001110001:ColourData=12'h2F2;
20'b00000100000001110001:ColourData=12'h4F2;
20'b00000100010001110001:ColourData=12'h3F1;
20'b00000100100001110001:ColourData=12'h3F1;
20'b00000100110001110001:ColourData=12'h6C0;
20'b00000101000001110001:ColourData=12'hB60;
20'b00000101010001110001:ColourData=12'hD30;
20'b00000101100001110001:ColourData=12'hD30;
20'b00000101110001110001:ColourData=12'hD30;
20'b00000110000001110001:ColourData=12'hE40;
20'b00000110010001110001:ColourData=12'hE40;
20'b00000110100001110001:ColourData=12'hE40;
20'b00000110110001110001:ColourData=12'hF40;
20'b00000111000001110001:ColourData=12'hE40;
20'b00000111010001110001:ColourData=12'h890;
20'b00000111100001110001:ColourData=12'h3F0;
20'b00000111110001110001:ColourData=12'h8F7;
20'b00000000000001110010:ColourData=12'h3F3;
20'b00000000010001110010:ColourData=12'h0F0;
20'b00000000100001110010:ColourData=12'h0F0;
20'b00000000110001110010:ColourData=12'h0F0;
20'b00000001000001110010:ColourData=12'h0F0;
20'b00000001010001110010:ColourData=12'h0F0;
20'b00000001100001110010:ColourData=12'h0F0;
20'b00000001110001110010:ColourData=12'h3F1;
20'b00000010000001110010:ColourData=12'h3F1;
20'b00000010010001110010:ColourData=12'h0F0;
20'b00000010100001110010:ColourData=12'h0F0;
20'b00000010110001110010:ColourData=12'h0F0;
20'b00000011000001110010:ColourData=12'h0F0;
20'b00000011010001110010:ColourData=12'h0F0;
20'b00000011100001110010:ColourData=12'h0F0;
20'b00000011110001110010:ColourData=12'h2F2;
20'b00000100000001110010:ColourData=12'h4F2;
20'b00000100010001110010:ColourData=12'h4F1;
20'b00000100100001110010:ColourData=12'h7C1;
20'b00000100110001110010:ColourData=12'hB70;
20'b00000101000001110010:ColourData=12'hA70;
20'b00000101010001110010:ColourData=12'hB70;
20'b00000101100001110010:ColourData=12'hB70;
20'b00000101110001110010:ColourData=12'hA70;
20'b00000110000001110010:ColourData=12'hC81;
20'b00000110010001110010:ColourData=12'hE82;
20'b00000110100001110010:ColourData=12'hC81;
20'b00000110110001110010:ColourData=12'hF93;
20'b00000111000001110010:ColourData=12'hCB3;
20'b00000111010001110010:ColourData=12'h6D1;
20'b00000111100001110010:ColourData=12'h4E1;
20'b00000111110001110010:ColourData=12'h8F7;
20'b00000000000001110011:ColourData=12'h3F3;
20'b00000000010001110011:ColourData=12'h0F0;
20'b00000000100001110011:ColourData=12'h0F0;
20'b00000000110001110011:ColourData=12'h0F0;
20'b00000001000001110011:ColourData=12'h0F0;
20'b00000001010001110011:ColourData=12'h0F0;
20'b00000001100001110011:ColourData=12'h0F0;
20'b00000001110001110011:ColourData=12'h3F1;
20'b00000010000001110011:ColourData=12'h3F1;
20'b00000010010001110011:ColourData=12'h0F0;
20'b00000010100001110011:ColourData=12'h0F0;
20'b00000010110001110011:ColourData=12'h0F0;
20'b00000011000001110011:ColourData=12'h0F0;
20'b00000011010001110011:ColourData=12'h0F0;
20'b00000011100001110011:ColourData=12'h0F0;
20'b00000011110001110011:ColourData=12'h2F2;
20'b00000100000001110011:ColourData=12'h4F2;
20'b00000100010001110011:ColourData=12'h6E1;
20'b00000100100001110011:ColourData=12'hF93;
20'b00000100110001110011:ColourData=12'hE82;
20'b00000101000001110011:ColourData=12'hB70;
20'b00000101010001110011:ColourData=12'hF93;
20'b00000101100001110011:ColourData=12'hD82;
20'b00000101110001110011:ColourData=12'hB70;
20'b00000110000001110011:ColourData=12'hE92;
20'b00000110010001110011:ColourData=12'hF93;
20'b00000110100001110011:ColourData=12'hE93;
20'b00000110110001110011:ColourData=12'hE82;
20'b00000111000001110011:ColourData=12'hE93;
20'b00000111010001110011:ColourData=12'hF93;
20'b00000111100001110011:ColourData=12'hBB2;
20'b00000111110001110011:ColourData=12'hAE7;
20'b00000000000001110100:ColourData=12'h3F3;
20'b00000000010001110100:ColourData=12'h0F0;
20'b00000000100001110100:ColourData=12'h0F0;
20'b00000000110001110100:ColourData=12'h0F0;
20'b00000001000001110100:ColourData=12'h0F0;
20'b00000001010001110100:ColourData=12'h0F0;
20'b00000001100001110100:ColourData=12'h0F0;
20'b00000001110001110100:ColourData=12'h3F1;
20'b00000010000001110100:ColourData=12'h3F1;
20'b00000010010001110100:ColourData=12'h0F0;
20'b00000010100001110100:ColourData=12'h0F0;
20'b00000010110001110100:ColourData=12'h0F0;
20'b00000011000001110100:ColourData=12'h0F0;
20'b00000011010001110100:ColourData=12'h0F0;
20'b00000011100001110100:ColourData=12'h0F0;
20'b00000011110001110100:ColourData=12'h2F2;
20'b00000100000001110100:ColourData=12'h4F2;
20'b00000100010001110100:ColourData=12'h5E1;
20'b00000100100001110100:ColourData=12'hDA3;
20'b00000100110001110100:ColourData=12'hE83;
20'b00000101000001110100:ColourData=12'hC81;
20'b00000101010001110100:ColourData=12'hE93;
20'b00000101100001110100:ColourData=12'hE93;
20'b00000101110001110100:ColourData=12'hB70;
20'b00000110000001110100:ColourData=12'hC81;
20'b00000110010001110100:ColourData=12'hF94;
20'b00000110100001110100:ColourData=12'hE92;
20'b00000110110001110100:ColourData=12'hA70;
20'b00000111000001110100:ColourData=12'hB70;
20'b00000111010001110100:ColourData=12'hE82;
20'b00000111100001110100:ColourData=12'hD92;
20'b00000111110001110100:ColourData=12'hDC8;
20'b00000000000001110101:ColourData=12'h3F3;
20'b00000000010001110101:ColourData=12'h0F0;
20'b00000000100001110101:ColourData=12'h0F0;
20'b00000000110001110101:ColourData=12'h0F0;
20'b00000001000001110101:ColourData=12'h0F0;
20'b00000001010001110101:ColourData=12'h0F0;
20'b00000001100001110101:ColourData=12'h0F0;
20'b00000001110001110101:ColourData=12'h3F1;
20'b00000010000001110101:ColourData=12'h3F1;
20'b00000010010001110101:ColourData=12'h0F0;
20'b00000010100001110101:ColourData=12'h0F0;
20'b00000010110001110101:ColourData=12'h0F0;
20'b00000011000001110101:ColourData=12'h0F0;
20'b00000011010001110101:ColourData=12'h0F0;
20'b00000011100001110101:ColourData=12'h0F0;
20'b00000011110001110101:ColourData=12'h2F2;
20'b00000100000001110101:ColourData=12'h4F2;
20'b00000100010001110101:ColourData=12'h3F1;
20'b00000100100001110101:ColourData=12'h5E1;
20'b00000100110001110101:ColourData=12'hDA3;
20'b00000101000001110101:ColourData=12'hE71;
20'b00000101010001110101:ColourData=12'hC60;
20'b00000101100001110101:ColourData=12'hE82;
20'b00000101110001110101:ColourData=12'hE82;
20'b00000110000001110101:ColourData=12'hE92;
20'b00000110010001110101:ColourData=12'hE82;
20'b00000110100001110101:ColourData=12'hF83;
20'b00000110110001110101:ColourData=12'hE92;
20'b00000111000001110101:ColourData=12'hB70;
20'b00000111010001110101:ColourData=12'hA80;
20'b00000111100001110101:ColourData=12'h6B0;
20'b00000111110001110101:ColourData=12'h8F7;
20'b00000000000001110110:ColourData=12'h3F3;
20'b00000000010001110110:ColourData=12'h0F0;
20'b00000000100001110110:ColourData=12'h0F0;
20'b00000000110001110110:ColourData=12'h0F0;
20'b00000001000001110110:ColourData=12'h0F0;
20'b00000001010001110110:ColourData=12'h0F0;
20'b00000001100001110110:ColourData=12'h0F0;
20'b00000001110001110110:ColourData=12'h3F1;
20'b00000010000001110110:ColourData=12'h3F1;
20'b00000010010001110110:ColourData=12'h0F0;
20'b00000010100001110110:ColourData=12'h0F0;
20'b00000010110001110110:ColourData=12'h0F0;
20'b00000011000001110110:ColourData=12'h0F0;
20'b00000011010001110110:ColourData=12'h0F0;
20'b00000011100001110110:ColourData=12'h0F0;
20'b00000011110001110110:ColourData=12'h2F2;
20'b00000100000001110110:ColourData=12'h4F2;
20'b00000100010001110110:ColourData=12'h3F1;
20'b00000100100001110110:ColourData=12'h4E1;
20'b00000100110001110110:ColourData=12'h8A0;
20'b00000101000001110110:ColourData=12'hF30;
20'b00000101010001110110:ColourData=12'hF40;
20'b00000101100001110110:ColourData=12'hE50;
20'b00000101110001110110:ColourData=12'hB70;
20'b00000110000001110110:ColourData=12'hA70;
20'b00000110010001110110:ColourData=12'hC40;
20'b00000110100001110110:ColourData=12'hE40;
20'b00000110110001110110:ColourData=12'hE92;
20'b00000111000001110110:ColourData=12'hE82;
20'b00000111010001110110:ColourData=12'hBA2;
20'b00000111100001110110:ColourData=12'h4E0;
20'b00000111110001110110:ColourData=12'h8F7;
20'b00000000000001110111:ColourData=12'h3F3;
20'b00000000010001110111:ColourData=12'h0F0;
20'b00000000100001110111:ColourData=12'h0F0;
20'b00000000110001110111:ColourData=12'h0F0;
20'b00000001000001110111:ColourData=12'h0F0;
20'b00000001010001110111:ColourData=12'h0F0;
20'b00000001100001110111:ColourData=12'h0F0;
20'b00000001110001110111:ColourData=12'h3F1;
20'b00000010000001110111:ColourData=12'h3F1;
20'b00000010010001110111:ColourData=12'h0F0;
20'b00000010100001110111:ColourData=12'h0F0;
20'b00000010110001110111:ColourData=12'h0F0;
20'b00000011000001110111:ColourData=12'h0F0;
20'b00000011010001110111:ColourData=12'h0F0;
20'b00000011100001110111:ColourData=12'h0F0;
20'b00000011110001110111:ColourData=12'h2F2;
20'b00000100000001110111:ColourData=12'h4F2;
20'b00000100010001110111:ColourData=12'h3F1;
20'b00000100100001110111:ColourData=12'h6C1;
20'b00000100110001110111:ColourData=12'hE30;
20'b00000101000001110111:ColourData=12'hE50;
20'b00000101010001110111:ColourData=12'hF93;
20'b00000101100001110111:ColourData=12'hF93;
20'b00000101110001110111:ColourData=12'hD82;
20'b00000110000001110111:ColourData=12'hB60;
20'b00000110010001110111:ColourData=12'hE30;
20'b00000110100001110111:ColourData=12'hC50;
20'b00000110110001110111:ColourData=12'hA70;
20'b00000111000001110111:ColourData=12'hA70;
20'b00000111010001110111:ColourData=12'hA70;
20'b00000111100001110111:ColourData=12'h7A0;
20'b00000111110001110111:ColourData=12'h8F7;
20'b00000000000001111000:ColourData=12'h3F3;
20'b00000000010001111000:ColourData=12'h0F0;
20'b00000000100001111000:ColourData=12'h0F0;
20'b00000000110001111000:ColourData=12'h0F0;
20'b00000001000001111000:ColourData=12'h0F0;
20'b00000001010001111000:ColourData=12'h0F0;
20'b00000001100001111000:ColourData=12'h0F0;
20'b00000001110001111000:ColourData=12'h3F1;
20'b00000010000001111000:ColourData=12'h3F1;
20'b00000010010001111000:ColourData=12'h0F0;
20'b00000010100001111000:ColourData=12'h0F0;
20'b00000010110001111000:ColourData=12'h0F0;
20'b00000011000001111000:ColourData=12'h0F0;
20'b00000011010001111000:ColourData=12'h0F0;
20'b00000011100001111000:ColourData=12'h0F0;
20'b00000011110001111000:ColourData=12'h2F2;
20'b00000100000001111000:ColourData=12'h4F2;
20'b00000100010001111000:ColourData=12'h3F1;
20'b00000100100001111000:ColourData=12'h6C1;
20'b00000100110001111000:ColourData=12'hE30;
20'b00000101000001111000:ColourData=12'hC60;
20'b00000101010001111000:ColourData=12'hF83;
20'b00000101100001111000:ColourData=12'hF94;
20'b00000101110001111000:ColourData=12'hD92;
20'b00000110000001111000:ColourData=12'hA70;
20'b00000110010001111000:ColourData=12'hA70;
20'b00000110100001111000:ColourData=12'hA70;
20'b00000110110001111000:ColourData=12'hA70;
20'b00000111000001111000:ColourData=12'hA70;
20'b00000111010001111000:ColourData=12'hA60;
20'b00000111100001111000:ColourData=12'h7A0;
20'b00000111110001111000:ColourData=12'h8F7;
20'b00000000000001111001:ColourData=12'h3F3;
20'b00000000010001111001:ColourData=12'h0F0;
20'b00000000100001111001:ColourData=12'h0F0;
20'b00000000110001111001:ColourData=12'h0F0;
20'b00000001000001111001:ColourData=12'h0F0;
20'b00000001010001111001:ColourData=12'h0F0;
20'b00000001100001111001:ColourData=12'h0F0;
20'b00000001110001111001:ColourData=12'h3F1;
20'b00000010000001111001:ColourData=12'h3F1;
20'b00000010010001111001:ColourData=12'h0F0;
20'b00000010100001111001:ColourData=12'h0F0;
20'b00000010110001111001:ColourData=12'h0F0;
20'b00000011000001111001:ColourData=12'h0F0;
20'b00000011010001111001:ColourData=12'h0F0;
20'b00000011100001111001:ColourData=12'h0F0;
20'b00000011110001111001:ColourData=12'h2F2;
20'b00000100000001111001:ColourData=12'h4F2;
20'b00000100010001111001:ColourData=12'h3F1;
20'b00000100100001111001:ColourData=12'h5D1;
20'b00000100110001111001:ColourData=12'hC50;
20'b00000101000001111001:ColourData=12'hF20;
20'b00000101010001111001:ColourData=12'hF40;
20'b00000101100001111001:ColourData=12'hF72;
20'b00000101110001111001:ColourData=12'hE71;
20'b00000110000001111001:ColourData=12'hA60;
20'b00000110010001111001:ColourData=12'hA70;
20'b00000110100001111001:ColourData=12'hA70;
20'b00000110110001111001:ColourData=12'hA70;
20'b00000111000001111001:ColourData=12'hA70;
20'b00000111010001111001:ColourData=12'hA70;
20'b00000111100001111001:ColourData=12'h6B0;
20'b00000111110001111001:ColourData=12'h8F7;
20'b00000000000001111010:ColourData=12'h3F3;
20'b00000000010001111010:ColourData=12'h0F0;
20'b00000000100001111010:ColourData=12'h0F0;
20'b00000000110001111010:ColourData=12'h0F0;
20'b00000001000001111010:ColourData=12'h0F0;
20'b00000001010001111010:ColourData=12'h0F0;
20'b00000001100001111010:ColourData=12'h0F0;
20'b00000001110001111010:ColourData=12'h3F1;
20'b00000010000001111010:ColourData=12'h3F1;
20'b00000010010001111010:ColourData=12'h0F0;
20'b00000010100001111010:ColourData=12'h0F0;
20'b00000010110001111010:ColourData=12'h0F0;
20'b00000011000001111010:ColourData=12'h0F0;
20'b00000011010001111010:ColourData=12'h0F0;
20'b00000011100001111010:ColourData=12'h0F0;
20'b00000011110001111010:ColourData=12'h2F2;
20'b00000100000001111010:ColourData=12'h4F2;
20'b00000100010001111010:ColourData=12'h3F1;
20'b00000100100001111010:ColourData=12'h3F1;
20'b00000100110001111010:ColourData=12'h6C1;
20'b00000101000001111010:ColourData=12'hE30;
20'b00000101010001111010:ColourData=12'hD30;
20'b00000101100001111010:ColourData=12'hD40;
20'b00000101110001111010:ColourData=12'hE30;
20'b00000110000001111010:ColourData=12'hD30;
20'b00000110010001111010:ColourData=12'hB60;
20'b00000110100001111010:ColourData=12'hB60;
20'b00000110110001111010:ColourData=12'hB60;
20'b00000111000001111010:ColourData=12'hA70;
20'b00000111010001111010:ColourData=12'h6B0;
20'b00000111100001111010:ColourData=12'h3F1;
20'b00000111110001111010:ColourData=12'h8F7;
20'b00000000000001111011:ColourData=12'h3F3;
20'b00000000010001111011:ColourData=12'h0F0;
20'b00000000100001111011:ColourData=12'h0F0;
20'b00000000110001111011:ColourData=12'h0F0;
20'b00000001000001111011:ColourData=12'h0F0;
20'b00000001010001111011:ColourData=12'h0F0;
20'b00000001100001111011:ColourData=12'h0F0;
20'b00000001110001111011:ColourData=12'h3F1;
20'b00000010000001111011:ColourData=12'h3F1;
20'b00000010010001111011:ColourData=12'h0F0;
20'b00000010100001111011:ColourData=12'h0F0;
20'b00000010110001111011:ColourData=12'h0F0;
20'b00000011000001111011:ColourData=12'h0F0;
20'b00000011010001111011:ColourData=12'h0F0;
20'b00000011100001111011:ColourData=12'h0F0;
20'b00000011110001111011:ColourData=12'h2F2;
20'b00000100000001111011:ColourData=12'h4F2;
20'b00000100010001111011:ColourData=12'h3F1;
20'b00000100100001111011:ColourData=12'h3F1;
20'b00000100110001111011:ColourData=12'h5D1;
20'b00000101000001111011:ColourData=12'hB60;
20'b00000101010001111011:ColourData=12'hA70;
20'b00000101100001111011:ColourData=12'hA70;
20'b00000101110001111011:ColourData=12'hB60;
20'b00000110000001111011:ColourData=12'hE30;
20'b00000110010001111011:ColourData=12'hF20;
20'b00000110100001111011:ColourData=12'hE30;
20'b00000110110001111011:ColourData=12'hF20;
20'b00000111000001111011:ColourData=12'hB70;
20'b00000111010001111011:ColourData=12'h3F1;
20'b00000111100001111011:ColourData=12'h3F0;
20'b00000111110001111011:ColourData=12'h8F7;
20'b00000000000001111100:ColourData=12'h3F3;
20'b00000000010001111100:ColourData=12'h0F0;
20'b00000000100001111100:ColourData=12'h0F0;
20'b00000000110001111100:ColourData=12'h0F0;
20'b00000001000001111100:ColourData=12'h0F0;
20'b00000001010001111100:ColourData=12'h0F0;
20'b00000001100001111100:ColourData=12'h0F0;
20'b00000001110001111100:ColourData=12'h3F1;
20'b00000010000001111100:ColourData=12'h3F1;
20'b00000010010001111100:ColourData=12'h0F0;
20'b00000010100001111100:ColourData=12'h0F0;
20'b00000010110001111100:ColourData=12'h0F0;
20'b00000011000001111100:ColourData=12'h0F0;
20'b00000011010001111100:ColourData=12'h0F0;
20'b00000011100001111100:ColourData=12'h0F0;
20'b00000011110001111100:ColourData=12'h2F2;
20'b00000100000001111100:ColourData=12'h4F2;
20'b00000100010001111100:ColourData=12'h4F1;
20'b00000100100001111100:ColourData=12'h5D1;
20'b00000100110001111100:ColourData=12'h5D1;
20'b00000101000001111100:ColourData=12'h6B0;
20'b00000101010001111100:ColourData=12'hB60;
20'b00000101100001111100:ColourData=12'hB60;
20'b00000101110001111100:ColourData=12'hA70;
20'b00000110000001111100:ColourData=12'hB60;
20'b00000110010001111100:ColourData=12'hE30;
20'b00000110100001111100:ColourData=12'hF20;
20'b00000110110001111100:ColourData=12'hE30;
20'b00000111000001111100:ColourData=12'h990;
20'b00000111010001111100:ColourData=12'h3F1;
20'b00000111100001111100:ColourData=12'h3F0;
20'b00000111110001111100:ColourData=12'h8F7;
20'b00000000000001111101:ColourData=12'h3F3;
20'b00000000010001111101:ColourData=12'h0F0;
20'b00000000100001111101:ColourData=12'h0F0;
20'b00000000110001111101:ColourData=12'h0F0;
20'b00000001000001111101:ColourData=12'h0F0;
20'b00000001010001111101:ColourData=12'h0F0;
20'b00000001100001111101:ColourData=12'h0F0;
20'b00000001110001111101:ColourData=12'h3F1;
20'b00000010000001111101:ColourData=12'h3F1;
20'b00000010010001111101:ColourData=12'h0F0;
20'b00000010100001111101:ColourData=12'h0F0;
20'b00000010110001111101:ColourData=12'h0F0;
20'b00000011000001111101:ColourData=12'h0F0;
20'b00000011010001111101:ColourData=12'h0F0;
20'b00000011100001111101:ColourData=12'h0F0;
20'b00000011110001111101:ColourData=12'h2F2;
20'b00000100000001111101:ColourData=12'h4F2;
20'b00000100010001111101:ColourData=12'h5D1;
20'b00000100100001111101:ColourData=12'hA70;
20'b00000100110001111101:ColourData=12'hA70;
20'b00000101000001111101:ColourData=12'hB60;
20'b00000101010001111101:ColourData=12'hD30;
20'b00000101100001111101:ColourData=12'hD40;
20'b00000101110001111101:ColourData=12'hB60;
20'b00000110000001111101:ColourData=12'hA70;
20'b00000110010001111101:ColourData=12'h980;
20'b00000110100001111101:ColourData=12'hC50;
20'b00000110110001111101:ColourData=12'h990;
20'b00000111000001111101:ColourData=12'h3F1;
20'b00000111010001111101:ColourData=12'h3F1;
20'b00000111100001111101:ColourData=12'h3F0;
20'b00000111110001111101:ColourData=12'h8F7;
20'b00000000000001111110:ColourData=12'h3F3;
20'b00000000010001111110:ColourData=12'h0F0;
20'b00000000100001111110:ColourData=12'h0F0;
20'b00000000110001111110:ColourData=12'h0F0;
20'b00000001000001111110:ColourData=12'h0F0;
20'b00000001010001111110:ColourData=12'h0F0;
20'b00000001100001111110:ColourData=12'h0F0;
20'b00000001110001111110:ColourData=12'h3F1;
20'b00000010000001111110:ColourData=12'h3F1;
20'b00000010010001111110:ColourData=12'h0F0;
20'b00000010100001111110:ColourData=12'h0F0;
20'b00000010110001111110:ColourData=12'h0F0;
20'b00000011000001111110:ColourData=12'h0F0;
20'b00000011010001111110:ColourData=12'h0F0;
20'b00000011100001111110:ColourData=12'h0F0;
20'b00000011110001111110:ColourData=12'h2F2;
20'b00000100000001111110:ColourData=12'h4F2;
20'b00000100010001111110:ColourData=12'h4E1;
20'b00000100100001111110:ColourData=12'h980;
20'b00000100110001111110:ColourData=12'hA70;
20'b00000101000001111110:ColourData=12'hA70;
20'b00000101010001111110:ColourData=12'hA70;
20'b00000101100001111110:ColourData=12'hB60;
20'b00000101110001111110:ColourData=12'hD40;
20'b00000110000001111110:ColourData=12'h980;
20'b00000110010001111110:ColourData=12'h3F1;
20'b00000110100001111110:ColourData=12'h3F1;
20'b00000110110001111110:ColourData=12'h3F1;
20'b00000111000001111110:ColourData=12'h3F1;
20'b00000111010001111110:ColourData=12'h3F1;
20'b00000111100001111110:ColourData=12'h3F0;
20'b00000111110001111110:ColourData=12'h8F7;
20'b00000000000001111111:ColourData=12'h3F3;
20'b00000000010001111111:ColourData=12'h0F0;
20'b00000000100001111111:ColourData=12'h0F0;
20'b00000000110001111111:ColourData=12'h0F0;
20'b00000001000001111111:ColourData=12'h0F0;
20'b00000001010001111111:ColourData=12'h0F0;
20'b00000001100001111111:ColourData=12'h0E0;
20'b00000001110001111111:ColourData=12'h2D1;
20'b00000010000001111111:ColourData=12'h3D1;
20'b00000010010001111111:ColourData=12'h0D0;
20'b00000010100001111111:ColourData=12'h0F0;
20'b00000010110001111111:ColourData=12'h0F0;
20'b00000011000001111111:ColourData=12'h0F0;
20'b00000011010001111111:ColourData=12'h0F0;
20'b00000011100001111111:ColourData=12'h0F0;
20'b00000011110001111111:ColourData=12'h2F2;
20'b00000100000001111111:ColourData=12'h4F2;
20'b00000100010001111111:ColourData=12'h3F1;
20'b00000100100001111111:ColourData=12'h4E1;
20'b00000100110001111111:ColourData=12'h890;
20'b00000101000001111111:ColourData=12'h890;
20'b00000101010001111111:ColourData=12'h890;
20'b00000101100001111111:ColourData=12'h890;
20'b00000101110001111111:ColourData=12'h7B0;
20'b00000110000001111111:ColourData=12'h3F1;
20'b00000110010001111111:ColourData=12'h3F1;
20'b00000110100001111111:ColourData=12'h3F1;
20'b00000110110001111111:ColourData=12'h3F1;
20'b00000111000001111111:ColourData=12'h4E1;
20'b00000111010001111111:ColourData=12'h6E1;
20'b00000111100001111111:ColourData=12'h6E1;
20'b00000111110001111111:ColourData=12'hAE7;
20'b00000000000010000000:ColourData=12'h3F3;
20'b00000000010010000000:ColourData=12'h0F0;
20'b00000000100010000000:ColourData=12'h0F0;
20'b00000000110010000000:ColourData=12'h0F0;
20'b00000001000010000000:ColourData=12'h0F0;
20'b00000001010010000000:ColourData=12'h0D0;
20'b00000001100010000000:ColourData=12'h040;
20'b00000001110010000000:ColourData=12'h010;
20'b00000010000010000000:ColourData=12'h010;
20'b00000010010010000000:ColourData=12'h020;
20'b00000010100010000000:ColourData=12'h0C0;
20'b00000010110010000000:ColourData=12'h0F0;
20'b00000011000010000000:ColourData=12'h0F0;
20'b00000011010010000000:ColourData=12'h0F0;
20'b00000011100010000000:ColourData=12'h0F0;
20'b00000011110010000000:ColourData=12'h2F2;
20'b00000100000010000000:ColourData=12'h4F2;
20'b00000100010010000000:ColourData=12'h3F1;
20'b00000100100010000000:ColourData=12'h3F1;
20'b00000100110010000000:ColourData=12'h3F1;
20'b00000101000010000000:ColourData=12'h3F1;
20'b00000101010010000000:ColourData=12'h4E1;
20'b00000101100010000000:ColourData=12'h6C1;
20'b00000101110010000000:ColourData=12'h6C1;
20'b00000110000010000000:ColourData=12'h6C1;
20'b00000110010010000000:ColourData=12'h6C1;
20'b00000110100010000000:ColourData=12'h6C1;
20'b00000110110010000000:ColourData=12'h5D1;
20'b00000111000010000000:ColourData=12'h7D2;
20'b00000111010010000000:ColourData=12'hF93;
20'b00000111100010000000:ColourData=12'hF93;
20'b00000111110010000000:ColourData=12'hFC8;
20'b00000000000010000001:ColourData=12'h3F3;
20'b00000000010010000001:ColourData=12'h0F0;
20'b00000000100010000001:ColourData=12'h0F0;
20'b00000000110010000001:ColourData=12'h0F0;
20'b00000001000010000001:ColourData=12'h0D0;
20'b00000001010010000001:ColourData=12'h040;
20'b00000001100010000001:ColourData=12'h2A0;
20'b00000001110010000001:ColourData=12'h170;
20'b00000010000010000001:ColourData=12'h160;
20'b00000010010010000001:ColourData=12'h160;
20'b00000010100010000001:ColourData=12'h030;
20'b00000010110010000001:ColourData=12'h0C0;
20'b00000011000010000001:ColourData=12'h0F0;
20'b00000011010010000001:ColourData=12'h0F0;
20'b00000011100010000001:ColourData=12'h0F0;
20'b00000011110010000001:ColourData=12'h2F2;
20'b00000100000010000001:ColourData=12'h4F2;
20'b00000100010010000001:ColourData=12'h3F1;
20'b00000100100010000001:ColourData=12'h3F1;
20'b00000100110010000001:ColourData=12'h3F1;
20'b00000101000010000001:ColourData=12'h4E1;
20'b00000101010010000001:ColourData=12'h8A0;
20'b00000101100010000001:ColourData=12'hF30;
20'b00000101110010000001:ColourData=12'hF20;
20'b00000110000010000001:ColourData=12'hE20;
20'b00000110010010000001:ColourData=12'hE20;
20'b00000110100010000001:ColourData=12'hF20;
20'b00000110110010000001:ColourData=12'hB60;
20'b00000111000010000001:ColourData=12'h9B1;
20'b00000111010010000001:ColourData=12'hF83;
20'b00000111100010000001:ColourData=12'hF93;
20'b00000111110010000001:ColourData=12'hFC8;
20'b00000000000010000010:ColourData=12'h3F3;
20'b00000000010010000010:ColourData=12'h0F0;
20'b00000000100010000010:ColourData=12'h0F0;
20'b00000000110010000010:ColourData=12'h0E0;
20'b00000001000010000010:ColourData=12'h040;
20'b00000001010010000010:ColourData=12'h2B1;
20'b00000001100010000010:ColourData=12'h290;
20'b00000001110010000010:ColourData=12'h170;
20'b00000010000010000010:ColourData=12'h170;
20'b00000010010010000010:ColourData=12'h170;
20'b00000010100010000010:ColourData=12'h160;
20'b00000010110010000010:ColourData=12'h020;
20'b00000011000010000010:ColourData=12'h0D0;
20'b00000011010010000010:ColourData=12'h0F0;
20'b00000011100010000010:ColourData=12'h0F0;
20'b00000011110010000010:ColourData=12'h2F2;
20'b00000100000010000010:ColourData=12'h4F2;
20'b00000100010010000010:ColourData=12'h3F1;
20'b00000100100010000010:ColourData=12'h3F1;
20'b00000100110010000010:ColourData=12'h3F1;
20'b00000101000010000010:ColourData=12'h6C1;
20'b00000101010010000010:ColourData=12'hD40;
20'b00000101100010000010:ColourData=12'hD30;
20'b00000101110010000010:ColourData=12'hE40;
20'b00000110000010000010:ColourData=12'hF40;
20'b00000110010010000010:ColourData=12'hE40;
20'b00000110100010000010:ColourData=12'hE40;
20'b00000110110010000010:ColourData=12'hF40;
20'b00000111000010000010:ColourData=12'hE40;
20'b00000111010010000010:ColourData=12'hE50;
20'b00000111100010000010:ColourData=12'hE92;
20'b00000111110010000010:ColourData=12'hEB8;
20'b00000000000010000011:ColourData=12'h3F3;
20'b00000000010010000011:ColourData=12'h0F0;
20'b00000000100010000011:ColourData=12'h0F0;
20'b00000000110010000011:ColourData=12'h0E0;
20'b00000001000010000011:ColourData=12'h020;
20'b00000001010010000011:ColourData=12'h2B1;
20'b00000001100010000011:ColourData=12'h280;
20'b00000001110010000011:ColourData=12'h170;
20'b00000010000010000011:ColourData=12'h170;
20'b00000010010010000011:ColourData=12'h170;
20'b00000010100010000011:ColourData=12'h160;
20'b00000010110010000011:ColourData=12'h010;
20'b00000011000010000011:ColourData=12'h0D0;
20'b00000011010010000011:ColourData=12'h0F0;
20'b00000011100010000011:ColourData=12'h0F0;
20'b00000011110010000011:ColourData=12'h2F2;
20'b00000100000010000011:ColourData=12'h4F2;
20'b00000100010010000011:ColourData=12'h3F1;
20'b00000100100010000011:ColourData=12'h3F1;
20'b00000100110010000011:ColourData=12'h4F1;
20'b00000101000010000011:ColourData=12'h6C0;
20'b00000101010010000011:ColourData=12'hB70;
20'b00000101100010000011:ColourData=12'hA70;
20'b00000101110010000011:ColourData=12'hC81;
20'b00000110000010000011:ColourData=12'hF93;
20'b00000110010010000011:ColourData=12'hD82;
20'b00000110100010000011:ColourData=12'hB70;
20'b00000110110010000011:ColourData=12'hF93;
20'b00000111000010000011:ColourData=12'hD82;
20'b00000111010010000011:ColourData=12'hA70;
20'b00000111100010000011:ColourData=12'hA60;
20'b00000111110010000011:ColourData=12'hCA6;
20'b00000000000010000100:ColourData=12'h3F3;
20'b00000000010010000100:ColourData=12'h0F0;
20'b00000000100010000100:ColourData=12'h0F0;
20'b00000000110010000100:ColourData=12'h0E0;
20'b00000001000010000100:ColourData=12'h020;
20'b00000001010010000100:ColourData=12'h160;
20'b00000001100010000100:ColourData=12'h170;
20'b00000001110010000100:ColourData=12'h170;
20'b00000010000010000100:ColourData=12'h170;
20'b00000010010010000100:ColourData=12'h170;
20'b00000010100010000100:ColourData=12'h160;
20'b00000010110010000100:ColourData=12'h010;
20'b00000011000010000100:ColourData=12'h0D0;
20'b00000011010010000100:ColourData=12'h0F0;
20'b00000011100010000100:ColourData=12'h0F0;
20'b00000011110010000100:ColourData=12'h2F2;
20'b00000100000010000100:ColourData=12'h4F2;
20'b00000100010010000100:ColourData=12'h3F1;
20'b00000100100010000100:ColourData=12'h3F1;
20'b00000100110010000100:ColourData=12'h5D0;
20'b00000101000010000100:ColourData=12'hB80;
20'b00000101010010000100:ColourData=12'hE92;
20'b00000101100010000100:ColourData=12'hB70;
20'b00000101110010000100:ColourData=12'hE92;
20'b00000110000010000100:ColourData=12'hF93;
20'b00000110010010000100:ColourData=12'hE92;
20'b00000110100010000100:ColourData=12'hC81;
20'b00000110110010000100:ColourData=12'hE93;
20'b00000111000010000100:ColourData=12'hE92;
20'b00000111010010000100:ColourData=12'hB70;
20'b00000111100010000100:ColourData=12'hA70;
20'b00000111110010000100:ColourData=12'hCA6;
20'b00000000000010000101:ColourData=12'h3F3;
20'b00000000010010000101:ColourData=12'h0F0;
20'b00000000100010000101:ColourData=12'h0F0;
20'b00000000110010000101:ColourData=12'h0E0;
20'b00000001000010000101:ColourData=12'h030;
20'b00000001010010000101:ColourData=12'h150;
20'b00000001100010000101:ColourData=12'h170;
20'b00000001110010000101:ColourData=12'h170;
20'b00000010000010000101:ColourData=12'h170;
20'b00000010010010000101:ColourData=12'h170;
20'b00000010100010000101:ColourData=12'h160;
20'b00000010110010000101:ColourData=12'h020;
20'b00000011000010000101:ColourData=12'h0D0;
20'b00000011010010000101:ColourData=12'h0F0;
20'b00000011100010000101:ColourData=12'h0F0;
20'b00000011110010000101:ColourData=12'h2F2;
20'b00000100000010000101:ColourData=12'h4F2;
20'b00000100010010000101:ColourData=12'h3F1;
20'b00000100100010000101:ColourData=12'h3F1;
20'b00000100110010000101:ColourData=12'h5D0;
20'b00000101000010000101:ColourData=12'hB70;
20'b00000101010010000101:ColourData=12'hD81;
20'b00000101100010000101:ColourData=12'hB70;
20'b00000101110010000101:ColourData=12'hC81;
20'b00000110000010000101:ColourData=12'hF93;
20'b00000110010010000101:ColourData=12'hF93;
20'b00000110100010000101:ColourData=12'hC81;
20'b00000110110010000101:ColourData=12'hB70;
20'b00000111000010000101:ColourData=12'hE92;
20'b00000111010010000101:ColourData=12'hE92;
20'b00000111100010000101:ColourData=12'hC80;
20'b00000111110010000101:ColourData=12'hCA6;
20'b00000000000010000110:ColourData=12'h3F3;
20'b00000000010010000110:ColourData=12'h0F0;
20'b00000000100010000110:ColourData=12'h0F0;
20'b00000000110010000110:ColourData=12'h0F0;
20'b00000001000010000110:ColourData=12'h0D0;
20'b00000001010010000110:ColourData=12'h030;
20'b00000001100010000110:ColourData=12'h150;
20'b00000001110010000110:ColourData=12'h160;
20'b00000010000010000110:ColourData=12'h160;
20'b00000010010010000110:ColourData=12'h160;
20'b00000010100010000110:ColourData=12'h030;
20'b00000010110010000110:ColourData=12'h0C0;
20'b00000011000010000110:ColourData=12'h0F0;
20'b00000011010010000110:ColourData=12'h0F0;
20'b00000011100010000110:ColourData=12'h0F0;
20'b00000011110010000110:ColourData=12'h2F2;
20'b00000100000010000110:ColourData=12'h4F2;
20'b00000100010010000110:ColourData=12'h3F1;
20'b00000100100010000110:ColourData=12'h3F1;
20'b00000100110010000110:ColourData=12'h4E1;
20'b00000101000010000110:ColourData=12'h890;
20'b00000101010010000110:ColourData=12'hA90;
20'b00000101100010000110:ColourData=12'hF93;
20'b00000101110010000110:ColourData=12'hF93;
20'b00000110000010000110:ColourData=12'hF93;
20'b00000110010010000110:ColourData=12'hE92;
20'b00000110100010000110:ColourData=12'hB70;
20'b00000110110010000110:ColourData=12'hB80;
20'b00000111000010000110:ColourData=12'hB70;
20'b00000111010010000110:ColourData=12'hA70;
20'b00000111100010000110:ColourData=12'h970;
20'b00000111110010000110:ColourData=12'hBB6;
20'b00000000000010000111:ColourData=12'h3F3;
20'b00000000010010000111:ColourData=12'h0F0;
20'b00000000100010000111:ColourData=12'h0F0;
20'b00000000110010000111:ColourData=12'h0F0;
20'b00000001000010000111:ColourData=12'h0F0;
20'b00000001010010000111:ColourData=12'h0D0;
20'b00000001100010000111:ColourData=12'h030;
20'b00000001110010000111:ColourData=12'h010;
20'b00000010000010000111:ColourData=12'h010;
20'b00000010010010000111:ColourData=12'h020;
20'b00000010100010000111:ColourData=12'h0C0;
20'b00000010110010000111:ColourData=12'h0F0;
20'b00000011000010000111:ColourData=12'h0F0;
20'b00000011010010000111:ColourData=12'h0F0;
20'b00000011100010000111:ColourData=12'h0F0;
20'b00000011110010000111:ColourData=12'h2F2;
20'b00000100000010000111:ColourData=12'h4F2;
20'b00000100010010000111:ColourData=12'h4F1;
20'b00000100100010000111:ColourData=12'h5D1;
20'b00000100110010000111:ColourData=12'h5D1;
20'b00000101000010000111:ColourData=12'h5D0;
20'b00000101010010000111:ColourData=12'h7C1;
20'b00000101100010000111:ColourData=12'hE82;
20'b00000101110010000111:ColourData=12'hF82;
20'b00000110000010000111:ColourData=12'hE92;
20'b00000110010010000111:ColourData=12'hE92;
20'b00000110100010000111:ColourData=12'hE82;
20'b00000110110010000111:ColourData=12'hF82;
20'b00000111000010000111:ColourData=12'hC81;
20'b00000111010010000111:ColourData=12'h970;
20'b00000111100010000111:ColourData=12'h6B0;
20'b00000111110010000111:ColourData=12'h8F7;
20'b00000000000010001000:ColourData=12'h3F3;
20'b00000000010010001000:ColourData=12'h0F0;
20'b00000000100010001000:ColourData=12'h0F0;
20'b00000000110010001000:ColourData=12'h0F0;
20'b00000001000010001000:ColourData=12'h0F0;
20'b00000001010010001000:ColourData=12'h0F0;
20'b00000001100010001000:ColourData=12'h0E0;
20'b00000001110010001000:ColourData=12'h2D1;
20'b00000010000010001000:ColourData=12'h3D1;
20'b00000010010010001000:ColourData=12'h0D0;
20'b00000010100010001000:ColourData=12'h0F0;
20'b00000010110010001000:ColourData=12'h0F0;
20'b00000011000010001000:ColourData=12'h0F0;
20'b00000011010010001000:ColourData=12'h0F0;
20'b00000011100010001000:ColourData=12'h0F0;
20'b00000011110010001000:ColourData=12'h2F2;
20'b00000100000010001000:ColourData=12'h4F2;
20'b00000100010010001000:ColourData=12'h6C0;
20'b00000100100010001000:ColourData=12'hA70;
20'b00000100110010001000:ColourData=12'hA70;
20'b00000101000010001000:ColourData=12'hA70;
20'b00000101010010001000:ColourData=12'hA70;
20'b00000101100010001000:ColourData=12'hB60;
20'b00000101110010001000:ColourData=12'hD40;
20'b00000110000010001000:ColourData=12'hB60;
20'b00000110010010001000:ColourData=12'hA70;
20'b00000110100010001000:ColourData=12'hB60;
20'b00000110110010001000:ColourData=12'hD40;
20'b00000111000010001000:ColourData=12'hB60;
20'b00000111010010001000:ColourData=12'h890;
20'b00000111100010001000:ColourData=12'h3E0;
20'b00000111110010001000:ColourData=12'h9E7;
20'b00000000000010001001:ColourData=12'h3F3;
20'b00000000010010001001:ColourData=12'h0F0;
20'b00000000100010001001:ColourData=12'h0F0;
20'b00000000110010001001:ColourData=12'h0F0;
20'b00000001000010001001:ColourData=12'h0F0;
20'b00000001010010001001:ColourData=12'h0F0;
20'b00000001100010001001:ColourData=12'h0F0;
20'b00000001110010001001:ColourData=12'h3F1;
20'b00000010000010001001:ColourData=12'h3F1;
20'b00000010010010001001:ColourData=12'h0F0;
20'b00000010100010001001:ColourData=12'h0F0;
20'b00000010110010001001:ColourData=12'h0F0;
20'b00000011000010001001:ColourData=12'h0F0;
20'b00000011010010001001:ColourData=12'h0F0;
20'b00000011100010001001:ColourData=12'h0F0;
20'b00000011110010001001:ColourData=12'h2F2;
20'b00000100000010001001:ColourData=12'h8D2;
20'b00000100010010001001:ColourData=12'hB70;
20'b00000100100010001001:ColourData=12'hA70;
20'b00000100110010001001:ColourData=12'hA70;
20'b00000101000010001001:ColourData=12'hA70;
20'b00000101010010001001:ColourData=12'hA70;
20'b00000101100010001001:ColourData=12'hA70;
20'b00000101110010001001:ColourData=12'hB60;
20'b00000110000010001001:ColourData=12'hD30;
20'b00000110010010001001:ColourData=12'hB60;
20'b00000110100010001001:ColourData=12'hB60;
20'b00000110110010001001:ColourData=12'hC50;
20'b00000111000010001001:ColourData=12'hF20;
20'b00000111010010001001:ColourData=12'hA80;
20'b00000111100010001001:ColourData=12'h5C0;
20'b00000111110010001001:ColourData=12'hCA6;
20'b00000000000010001010:ColourData=12'h3F3;
20'b00000000010010001010:ColourData=12'h0F0;
20'b00000000100010001010:ColourData=12'h0F0;
20'b00000000110010001010:ColourData=12'h0F0;
20'b00000001000010001010:ColourData=12'h0F0;
20'b00000001010010001010:ColourData=12'h0F0;
20'b00000001100010001010:ColourData=12'h0F0;
20'b00000001110010001010:ColourData=12'h3F1;
20'b00000010000010001010:ColourData=12'h3F1;
20'b00000010010010001010:ColourData=12'h0F0;
20'b00000010100010001010:ColourData=12'h0F0;
20'b00000010110010001010:ColourData=12'h0F0;
20'b00000011000010001010:ColourData=12'h0F0;
20'b00000011010010001010:ColourData=12'h0F0;
20'b00000011100010001010:ColourData=12'h0F0;
20'b00000011110010001010:ColourData=12'h3E2;
20'b00000100000010001010:ColourData=12'hFA4;
20'b00000100010010001010:ColourData=12'hE92;
20'b00000100100010001010:ColourData=12'hB70;
20'b00000100110010001010:ColourData=12'hB70;
20'b00000101000010001010:ColourData=12'hB60;
20'b00000101010010001010:ColourData=12'hB60;
20'b00000101100010001010:ColourData=12'hA70;
20'b00000101110010001010:ColourData=12'hC50;
20'b00000110000010001010:ColourData=12'hF30;
20'b00000110010010001010:ColourData=12'hF40;
20'b00000110100010001010:ColourData=12'hE20;
20'b00000110110010001010:ColourData=12'hF30;
20'b00000111000010001010:ColourData=12'hF30;
20'b00000111010010001010:ColourData=12'hB70;
20'b00000111100010001010:ColourData=12'h6B0;
20'b00000111110010001010:ColourData=12'hCA6;
20'b00000000000010001011:ColourData=12'h3F3;
20'b00000000010010001011:ColourData=12'h0F0;
20'b00000000100010001011:ColourData=12'h0F0;
20'b00000000110010001011:ColourData=12'h0F0;
20'b00000001000010001011:ColourData=12'h0F0;
20'b00000001010010001011:ColourData=12'h0F0;
20'b00000001100010001011:ColourData=12'h0F0;
20'b00000001110010001011:ColourData=12'h3F1;
20'b00000010000010001011:ColourData=12'h3F1;
20'b00000010010010001011:ColourData=12'h0F0;
20'b00000010100010001011:ColourData=12'h0F0;
20'b00000010110010001011:ColourData=12'h0F0;
20'b00000011000010001011:ColourData=12'h0F0;
20'b00000011010010001011:ColourData=12'h0F0;
20'b00000011100010001011:ColourData=12'h0F0;
20'b00000011110010001011:ColourData=12'h3E2;
20'b00000100000010001011:ColourData=12'hDB3;
20'b00000100010010001011:ColourData=12'hF93;
20'b00000100100010001011:ColourData=12'hF93;
20'b00000100110010001011:ColourData=12'hE71;
20'b00000101000010001011:ColourData=12'hF20;
20'b00000101010010001011:ColourData=12'hD30;
20'b00000101100010001011:ColourData=12'hC50;
20'b00000101110010001011:ColourData=12'hE20;
20'b00000110000010001011:ColourData=12'hF40;
20'b00000110010010001011:ColourData=12'hF61;
20'b00000110100010001011:ColourData=12'hF20;
20'b00000110110010001011:ColourData=12'hF40;
20'b00000111000010001011:ColourData=12'hF61;
20'b00000111010010001011:ColourData=12'hD40;
20'b00000111100010001011:ColourData=12'h970;
20'b00000111110010001011:ColourData=12'hCA6;
20'b00000000000010001100:ColourData=12'h3F3;
20'b00000000010010001100:ColourData=12'h0F0;
20'b00000000100010001100:ColourData=12'h0F0;
20'b00000000110010001100:ColourData=12'h0F0;
20'b00000001000010001100:ColourData=12'h0F0;
20'b00000001010010001100:ColourData=12'h0F0;
20'b00000001100010001100:ColourData=12'h0F0;
20'b00000001110010001100:ColourData=12'h3F1;
20'b00000010000010001100:ColourData=12'h3F1;
20'b00000010010010001100:ColourData=12'h0F0;
20'b00000010100010001100:ColourData=12'h0F0;
20'b00000010110010001100:ColourData=12'h0F0;
20'b00000011000010001100:ColourData=12'h0F0;
20'b00000011010010001100:ColourData=12'h0F0;
20'b00000011100010001100:ColourData=12'h0F0;
20'b00000011110010001100:ColourData=12'h2F2;
20'b00000100000010001100:ColourData=12'h6E2;
20'b00000100010010001100:ColourData=12'hCB2;
20'b00000100100010001100:ColourData=12'hD81;
20'b00000100110010001100:ColourData=12'hB60;
20'b00000101000010001100:ColourData=12'hE30;
20'b00000101010010001100:ColourData=12'hF30;
20'b00000101100010001100:ColourData=12'hF30;
20'b00000101110010001100:ColourData=12'hF30;
20'b00000110000010001100:ColourData=12'hF30;
20'b00000110010010001100:ColourData=12'hF30;
20'b00000110100010001100:ColourData=12'hF30;
20'b00000110110010001100:ColourData=12'hF20;
20'b00000111000010001100:ColourData=12'hF20;
20'b00000111010010001100:ColourData=12'hD40;
20'b00000111100010001100:ColourData=12'hA60;
20'b00000111110010001100:ColourData=12'hCA6;
20'b00000000000010001101:ColourData=12'h3F3;
20'b00000000010010001101:ColourData=12'h0F0;
20'b00000000100010001101:ColourData=12'h0F0;
20'b00000000110010001101:ColourData=12'h0F0;
20'b00000001000010001101:ColourData=12'h0F0;
20'b00000001010010001101:ColourData=12'h0F0;
20'b00000001100010001101:ColourData=12'h0F0;
20'b00000001110010001101:ColourData=12'h3F1;
20'b00000010000010001101:ColourData=12'h3F1;
20'b00000010010010001101:ColourData=12'h0F0;
20'b00000010100010001101:ColourData=12'h0F0;
20'b00000010110010001101:ColourData=12'h0F0;
20'b00000011000010001101:ColourData=12'h0F0;
20'b00000011010010001101:ColourData=12'h0F0;
20'b00000011100010001101:ColourData=12'h0F0;
20'b00000011110010001101:ColourData=12'h2F2;
20'b00000100000010001101:ColourData=12'h4F2;
20'b00000100010010001101:ColourData=12'h6C0;
20'b00000100100010001101:ColourData=12'hA70;
20'b00000100110010001101:ColourData=12'hA60;
20'b00000101000010001101:ColourData=12'hC50;
20'b00000101010010001101:ColourData=12'hF30;
20'b00000101100010001101:ColourData=12'hF30;
20'b00000101110010001101:ColourData=12'hF30;
20'b00000110000010001101:ColourData=12'hF20;
20'b00000110010010001101:ColourData=12'hF20;
20'b00000110100010001101:ColourData=12'hF20;
20'b00000110110010001101:ColourData=12'hE30;
20'b00000111000010001101:ColourData=12'hC50;
20'b00000111010010001101:ColourData=12'hB70;
20'b00000111100010001101:ColourData=12'h890;
20'b00000111110010001101:ColourData=12'hBB6;
20'b00000000000010001110:ColourData=12'h2F2;
20'b00000000010010001110:ColourData=12'h0F0;
20'b00000000100010001110:ColourData=12'h0F0;
20'b00000000110010001110:ColourData=12'h0F0;
20'b00000001000010001110:ColourData=12'h0F0;
20'b00000001010010001110:ColourData=12'h0F0;
20'b00000001100010001110:ColourData=12'h0F0;
20'b00000001110010001110:ColourData=12'h3F1;
20'b00000010000010001110:ColourData=12'h3F1;
20'b00000010010010001110:ColourData=12'h0F0;
20'b00000010100010001110:ColourData=12'h0F0;
20'b00000010110010001110:ColourData=12'h0F0;
20'b00000011000010001110:ColourData=12'h0F0;
20'b00000011010010001110:ColourData=12'h0F0;
20'b00000011100010001110:ColourData=12'h0F0;
20'b00000011110010001110:ColourData=12'h2F2;
20'b00000100000010001110:ColourData=12'h5D1;
20'b00000100010010001110:ColourData=12'hA70;
20'b00000100100010001110:ColourData=12'h970;
20'b00000100110010001110:ColourData=12'hA70;
20'b00000101000010001110:ColourData=12'hF20;
20'b00000101010010001110:ColourData=12'hF20;
20'b00000101100010001110:ColourData=12'hF20;
20'b00000101110010001110:ColourData=12'hF20;
20'b00000110000010001110:ColourData=12'hE30;
20'b00000110010010001110:ColourData=12'hC50;
20'b00000110100010001110:ColourData=12'hC50;
20'b00000110110010001110:ColourData=12'h990;
20'b00000111000010001110:ColourData=12'h3F1;
20'b00000111010010001110:ColourData=12'h3F1;
20'b00000111100010001110:ColourData=12'h3F0;
20'b00000111110010001110:ColourData=12'h8F7;
20'b00000000000010001111:ColourData=12'h3E4;
20'b00000000010010001111:ColourData=12'h0E0;
20'b00000000100010001111:ColourData=12'h0E0;
20'b00000000110010001111:ColourData=12'h0E0;
20'b00000001000010001111:ColourData=12'h0E0;
20'b00000001010010001111:ColourData=12'h0E0;
20'b00000001100010001111:ColourData=12'h0E0;
20'b00000001110010001111:ColourData=12'h4E1;
20'b00000010000010001111:ColourData=12'h4E1;
20'b00000010010010001111:ColourData=12'h1E0;
20'b00000010100010001111:ColourData=12'h0E0;
20'b00000010110010001111:ColourData=12'h0E0;
20'b00000011000010001111:ColourData=12'h0E0;
20'b00000011010010001111:ColourData=12'h0E0;
20'b00000011100010001111:ColourData=12'h0E0;
20'b00000011110010001111:ColourData=12'h2F3;
20'b00000100000010001111:ColourData=12'h5E2;
20'b00000100010010001111:ColourData=12'h890;
20'b00000100100010001111:ColourData=12'h7A0;
20'b00000100110010001111:ColourData=12'h5D1;
20'b00000101000010001111:ColourData=12'hC60;
20'b00000101010010001111:ColourData=12'hC60;
20'b00000101100010001111:ColourData=12'hC60;
20'b00000101110010001111:ColourData=12'hC50;
20'b00000110000010001111:ColourData=12'h990;
20'b00000110010010001111:ColourData=12'h3F1;
20'b00000110100010001111:ColourData=12'h3F1;
20'b00000110110010001111:ColourData=12'h3F1;
20'b00000111000010001111:ColourData=12'h3F1;
20'b00000111010010001111:ColourData=12'h3F1;
20'b00000111100010001111:ColourData=12'h3F0;
20'b00000111110010001111:ColourData=12'h8F7;
20'b00000000000010010000:ColourData=12'h8AC;
20'b00000000010010010000:ColourData=12'h963;
20'b00000000100010010000:ColourData=12'hA51;
20'b00000000110010010000:ColourData=12'hA51;
20'b00000001000010010000:ColourData=12'hA51;
20'b00000001010010010000:ColourData=12'hA51;
20'b00000001100010010000:ColourData=12'hA51;
20'b00000001110010010000:ColourData=12'hA51;
20'b00000010000010010000:ColourData=12'hB51;
20'b00000010010010010000:ColourData=12'hA51;
20'b00000010100010010000:ColourData=12'hA51;
20'b00000010110010010000:ColourData=12'hA51;
20'b00000011000010010000:ColourData=12'hA51;
20'b00000011010010010000:ColourData=12'hA51;
20'b00000011100010010000:ColourData=12'h952;
20'b00000011110010010000:ColourData=12'h6AA;
20'b00000100000010010000:ColourData=12'h4F2;
20'b00000100010010010000:ColourData=12'h3F1;
20'b00000100100010010000:ColourData=12'h3F1;
20'b00000100110010010000:ColourData=12'h4F1;
20'b00000101000010010000:ColourData=12'h6C1;
20'b00000101010010010000:ColourData=12'h6C1;
20'b00000101100010010000:ColourData=12'h6C1;
20'b00000101110010010000:ColourData=12'h6C1;
20'b00000110000010010000:ColourData=12'h6C1;
20'b00000110010010010000:ColourData=12'h5D1;
20'b00000110100010010000:ColourData=12'h3F1;
20'b00000110110010010000:ColourData=12'h3F1;
20'b00000111000010010000:ColourData=12'h3F1;
20'b00000111010010010000:ColourData=12'h3F1;
20'b00000111100010010000:ColourData=12'h3F0;
20'b00000111110010010000:ColourData=12'h8F7;
20'b00000000000010010001:ColourData=12'hC65;
20'b00000000010010010001:ColourData=12'hD72;
20'b00000000100010010001:ColourData=12'hD73;
20'b00000000110010010001:ColourData=12'hE83;
20'b00000001000010010001:ColourData=12'hE83;
20'b00000001010010010001:ColourData=12'hE83;
20'b00000001100010010001:ColourData=12'hE83;
20'b00000001110010010001:ColourData=12'hE83;
20'b00000010000010010001:ColourData=12'hE83;
20'b00000010010010010001:ColourData=12'hE83;
20'b00000010100010010001:ColourData=12'hE83;
20'b00000010110010010001:ColourData=12'hE83;
20'b00000011000010010001:ColourData=12'hE83;
20'b00000011010010010001:ColourData=12'hD73;
20'b00000011100010010001:ColourData=12'hC62;
20'b00000011110010010001:ColourData=12'h453;
20'b00000100000010010001:ColourData=12'h4F2;
20'b00000100010010010001:ColourData=12'h3F1;
20'b00000100100010010001:ColourData=12'h4E1;
20'b00000100110010010001:ColourData=12'h8A0;
20'b00000101000010010001:ColourData=12'hE30;
20'b00000101010010010001:ColourData=12'hF30;
20'b00000101100010010001:ColourData=12'hE30;
20'b00000101110010010001:ColourData=12'hE30;
20'b00000110000010010001:ColourData=12'hF20;
20'b00000110010010010001:ColourData=12'hC50;
20'b00000110100010010001:ColourData=12'h6C0;
20'b00000110110010010001:ColourData=12'h6C1;
20'b00000111000010010001:ColourData=12'h5D1;
20'b00000111010010010001:ColourData=12'h3F1;
20'b00000111100010010001:ColourData=12'h3F0;
20'b00000111110010010001:ColourData=12'h8F7;
20'b00000000000010010010:ColourData=12'hC64;
20'b00000000010010010010:ColourData=12'hD72;
20'b00000000100010010010:ColourData=12'h531;
20'b00000000110010010010:ColourData=12'hC72;
20'b00000001000010010010:ColourData=12'hF93;
20'b00000001010010010010:ColourData=12'hE83;
20'b00000001100010010010:ColourData=12'hE83;
20'b00000001110010010010:ColourData=12'hE83;
20'b00000010000010010010:ColourData=12'hE83;
20'b00000010010010010010:ColourData=12'hE83;
20'b00000010100010010010:ColourData=12'hE93;
20'b00000010110010010010:ColourData=12'hF93;
20'b00000011000010010010:ColourData=12'hD83;
20'b00000011010010010010:ColourData=12'h531;
20'b00000011100010010010:ColourData=12'hB62;
20'b00000011110010010010:ColourData=12'h342;
20'b00000100000010010010:ColourData=12'h4F2;
20'b00000100010010010010:ColourData=12'h3F1;
20'b00000100100010010010:ColourData=12'h5D1;
20'b00000100110010010010:ColourData=12'hD40;
20'b00000101000010010010:ColourData=12'hD30;
20'b00000101010010010010:ColourData=12'hE40;
20'b00000101100010010010:ColourData=12'hF40;
20'b00000101110010010010:ColourData=12'hE40;
20'b00000110000010010010:ColourData=12'hE40;
20'b00000110010010010010:ColourData=12'hF40;
20'b00000110100010010010:ColourData=12'hE50;
20'b00000110110010010010:ColourData=12'hC50;
20'b00000111000010010010:ColourData=12'h990;
20'b00000111010010010010:ColourData=12'h3F1;
20'b00000111100010010010:ColourData=12'h3F0;
20'b00000111110010010010:ColourData=12'h8F7;
20'b00000000000010010011:ColourData=12'hC64;
20'b00000000010010010011:ColourData=12'hD72;
20'b00000000100010010011:ColourData=12'hD83;
20'b00000000110010010011:ColourData=12'hE83;
20'b00000001000010010011:ColourData=12'hE83;
20'b00000001010010010011:ColourData=12'hC51;
20'b00000001100010010011:ColourData=12'hA41;
20'b00000001110010010011:ColourData=12'hA41;
20'b00000010000010010011:ColourData=12'hA41;
20'b00000010010010010011:ColourData=12'hB41;
20'b00000010100010010011:ColourData=12'hE83;
20'b00000010110010010011:ColourData=12'hE93;
20'b00000011000010010011:ColourData=12'hE83;
20'b00000011010010010011:ColourData=12'hD83;
20'b00000011100010010011:ColourData=12'hC72;
20'b00000011110010010011:ColourData=12'h342;
20'b00000100000010010011:ColourData=12'h4F2;
20'b00000100010010010011:ColourData=12'h3F1;
20'b00000100100010010011:ColourData=12'h6C0;
20'b00000100110010010011:ColourData=12'hB70;
20'b00000101000010010011:ColourData=12'hA70;
20'b00000101010010010011:ColourData=12'hC81;
20'b00000101100010010011:ColourData=12'hF93;
20'b00000101110010010011:ColourData=12'hD82;
20'b00000110000010010011:ColourData=12'hB70;
20'b00000110010010010011:ColourData=12'hF93;
20'b00000110100010010011:ColourData=12'hCA3;
20'b00000110110010010011:ColourData=12'h6D1;
20'b00000111000010010011:ColourData=12'h5E1;
20'b00000111010010010011:ColourData=12'h3F1;
20'b00000111100010010011:ColourData=12'h3F0;
20'b00000111110010010011:ColourData=12'h8F7;
20'b00000000000010010100:ColourData=12'hC64;
20'b00000000010010010100:ColourData=12'hD72;
20'b00000000100010010100:ColourData=12'hF93;
20'b00000000110010010100:ColourData=12'hE83;
20'b00000001000010010100:ColourData=12'hC51;
20'b00000001010010010100:ColourData=12'hA31;
20'b00000001100010010100:ColourData=12'h200;
20'b00000001110010010100:ColourData=12'h100;
20'b00000010000010010100:ColourData=12'h210;
20'b00000010010010010100:ColourData=12'hA31;
20'b00000010100010010100:ColourData=12'hC41;
20'b00000010110010010100:ColourData=12'hD73;
20'b00000011000010010100:ColourData=12'hE83;
20'b00000011010010010100:ColourData=12'hF93;
20'b00000011100010010100:ColourData=12'hC72;
20'b00000011110010010100:ColourData=12'h342;
20'b00000100000010010100:ColourData=12'h4F2;
20'b00000100010010010100:ColourData=12'h5D0;
20'b00000100100010010100:ColourData=12'hB80;
20'b00000100110010010100:ColourData=12'hE82;
20'b00000101000010010100:ColourData=12'hB70;
20'b00000101010010010100:ColourData=12'hE92;
20'b00000101100010010100:ColourData=12'hF93;
20'b00000101110010010100:ColourData=12'hE92;
20'b00000110000010010100:ColourData=12'hC81;
20'b00000110010010010100:ColourData=12'hE93;
20'b00000110100010010100:ColourData=12'hF93;
20'b00000110110010010100:ColourData=12'hF93;
20'b00000111000010010100:ColourData=12'hCB3;
20'b00000111010010010100:ColourData=12'h5E1;
20'b00000111100010010100:ColourData=12'h3F0;
20'b00000111110010010100:ColourData=12'h8F7;
20'b00000000000010010101:ColourData=12'hC64;
20'b00000000010010010101:ColourData=12'hD72;
20'b00000000100010010101:ColourData=12'hE93;
20'b00000000110010010101:ColourData=12'hE83;
20'b00000001000010010101:ColourData=12'hC41;
20'b00000001010010010101:ColourData=12'hA31;
20'b00000001100010010101:ColourData=12'h100;
20'b00000001110010010101:ColourData=12'hA62;
20'b00000010000010010101:ColourData=12'hD73;
20'b00000010010010010101:ColourData=12'hB41;
20'b00000010100010010101:ColourData=12'hA31;
20'b00000010110010010101:ColourData=12'h310;
20'b00000011000010010101:ColourData=12'hD83;
20'b00000011010010010101:ColourData=12'hF93;
20'b00000011100010010101:ColourData=12'hC72;
20'b00000011110010010101:ColourData=12'h342;
20'b00000100000010010101:ColourData=12'h4F2;
20'b00000100010010010101:ColourData=12'h5D0;
20'b00000100100010010101:ColourData=12'hB70;
20'b00000100110010010101:ColourData=12'hD82;
20'b00000101000010010101:ColourData=12'hB70;
20'b00000101010010010101:ColourData=12'hC81;
20'b00000101100010010101:ColourData=12'hF93;
20'b00000101110010010101:ColourData=12'hF93;
20'b00000110000010010101:ColourData=12'hC81;
20'b00000110010010010101:ColourData=12'hB70;
20'b00000110100010010101:ColourData=12'hE82;
20'b00000110110010010101:ColourData=12'hE82;
20'b00000111000010010101:ColourData=12'hD92;
20'b00000111010010010101:ColourData=12'h9C2;
20'b00000111100010010101:ColourData=12'h3F0;
20'b00000111110010010101:ColourData=12'h8F7;
20'b00000000000010010110:ColourData=12'hC64;
20'b00000000010010010110:ColourData=12'hD72;
20'b00000000100010010110:ColourData=12'hE93;
20'b00000000110010010110:ColourData=12'hE83;
20'b00000001000010010110:ColourData=12'hC51;
20'b00000001010010010110:ColourData=12'h931;
20'b00000001100010010110:ColourData=12'h100;
20'b00000001110010010110:ColourData=12'hC73;
20'b00000010000010010110:ColourData=12'hE83;
20'b00000010010010010110:ColourData=12'hC41;
20'b00000010100010010110:ColourData=12'hA31;
20'b00000010110010010110:ColourData=12'h200;
20'b00000011000010010110:ColourData=12'hD73;
20'b00000011010010010110:ColourData=12'hF93;
20'b00000011100010010110:ColourData=12'hC72;
20'b00000011110010010110:ColourData=12'h342;
20'b00000100000010010110:ColourData=12'h4F2;
20'b00000100010010010110:ColourData=12'h4E1;
20'b00000100100010010110:ColourData=12'h890;
20'b00000100110010010110:ColourData=12'hA90;
20'b00000101000010010110:ColourData=12'hF93;
20'b00000101010010010110:ColourData=12'hF93;
20'b00000101100010010110:ColourData=12'hF94;
20'b00000101110010010110:ColourData=12'hE93;
20'b00000110000010010110:ColourData=12'hB70;
20'b00000110010010010110:ColourData=12'hB70;
20'b00000110100010010110:ColourData=12'hB70;
20'b00000110110010010110:ColourData=12'hA80;
20'b00000111000010010110:ColourData=12'h6B0;
20'b00000111010010010110:ColourData=12'h3F1;
20'b00000111100010010110:ColourData=12'h3F0;
20'b00000111110010010110:ColourData=12'h8F7;
20'b00000000000010010111:ColourData=12'hC64;
20'b00000000010010010111:ColourData=12'hD72;
20'b00000000100010010111:ColourData=12'hE93;
20'b00000000110010010111:ColourData=12'hE93;
20'b00000001000010010111:ColourData=12'hE83;
20'b00000001010010010111:ColourData=12'h420;
20'b00000001100010010111:ColourData=12'h100;
20'b00000001110010010111:ColourData=12'hC72;
20'b00000010000010010111:ColourData=12'hC51;
20'b00000010010010010111:ColourData=12'hA31;
20'b00000010100010010111:ColourData=12'h830;
20'b00000010110010010111:ColourData=12'h100;
20'b00000011000010010111:ColourData=12'hD73;
20'b00000011010010010111:ColourData=12'hF93;
20'b00000011100010010111:ColourData=12'hC72;
20'b00000011110010010111:ColourData=12'h342;
20'b00000100000010010111:ColourData=12'h4F2;
20'b00000100010010010111:ColourData=12'h3F1;
20'b00000100100010010111:ColourData=12'h3F1;
20'b00000100110010010111:ColourData=12'h6D1;
20'b00000101000010010111:ColourData=12'hF72;
20'b00000101010010010111:ColourData=12'hF72;
20'b00000101100010010111:ColourData=12'hE82;
20'b00000101110010010111:ColourData=12'hE82;
20'b00000110000010010111:ColourData=12'hD82;
20'b00000110010010010111:ColourData=12'hD82;
20'b00000110100010010111:ColourData=12'hE82;
20'b00000110110010010111:ColourData=12'hCA3;
20'b00000111000010010111:ColourData=12'h6D2;
20'b00000111010010010111:ColourData=12'h5E1;
20'b00000111100010010111:ColourData=12'h3F0;
20'b00000111110010010111:ColourData=12'h8F7;
20'b00000000000010011000:ColourData=12'hC64;
20'b00000000010010011000:ColourData=12'hD72;
20'b00000000100010011000:ColourData=12'hE93;
20'b00000000110010011000:ColourData=12'hE83;
20'b00000001000010011000:ColourData=12'hE93;
20'b00000001010010011000:ColourData=12'hE83;
20'b00000001100010011000:ColourData=12'hD83;
20'b00000001110010011000:ColourData=12'hC51;
20'b00000010000010011000:ColourData=12'hA31;
20'b00000010010010011000:ColourData=12'h100;
20'b00000010100010011000:ColourData=12'h100;
20'b00000010110010011000:ColourData=12'h210;
20'b00000011000010011000:ColourData=12'hD83;
20'b00000011010010011000:ColourData=12'hF93;
20'b00000011100010011000:ColourData=12'hC72;
20'b00000011110010011000:ColourData=12'h342;
20'b00000100000010011000:ColourData=12'h4F2;
20'b00000100010010011000:ColourData=12'h3F1;
20'b00000100100010011000:ColourData=12'h3F1;
20'b00000100110010011000:ColourData=12'h8A0;
20'b00000101000010011000:ColourData=12'hE30;
20'b00000101010010011000:ColourData=12'hC40;
20'b00000101100010011000:ColourData=12'hA70;
20'b00000101110010011000:ColourData=12'hA70;
20'b00000110000010011000:ColourData=12'hA70;
20'b00000110010010011000:ColourData=12'hA70;
20'b00000110100010011000:ColourData=12'hB70;
20'b00000110110010011000:ColourData=12'hF93;
20'b00000111000010011000:ColourData=12'hF93;
20'b00000111010010011000:ColourData=12'hCB3;
20'b00000111100010011000:ColourData=12'h4E1;
20'b00000111110010011000:ColourData=12'h8F7;
20'b00000000000010011001:ColourData=12'hC64;
20'b00000000010010011001:ColourData=12'hD72;
20'b00000000100010011001:ColourData=12'hE93;
20'b00000000110010011001:ColourData=12'hE83;
20'b00000001000010011001:ColourData=12'hE83;
20'b00000001010010011001:ColourData=12'hE93;
20'b00000001100010011001:ColourData=12'hE83;
20'b00000001110010011001:ColourData=12'hC51;
20'b00000010000010011001:ColourData=12'h931;
20'b00000010010010011001:ColourData=12'h100;
20'b00000010100010011001:ColourData=12'hB62;
20'b00000010110010011001:ColourData=12'hD83;
20'b00000011000010011001:ColourData=12'hE83;
20'b00000011010010011001:ColourData=12'hF93;
20'b00000011100010011001:ColourData=12'hC72;
20'b00000011110010011001:ColourData=12'h342;
20'b00000100000010011001:ColourData=12'h4F2;
20'b00000100010010011001:ColourData=12'h4E1;
20'b00000100100010011001:ColourData=12'h8A0;
20'b00000100110010011001:ColourData=12'hE30;
20'b00000101000010011001:ColourData=12'hD40;
20'b00000101010010011001:ColourData=12'hA70;
20'b00000101100010011001:ColourData=12'hA70;
20'b00000101110010011001:ColourData=12'hA70;
20'b00000110000010011001:ColourData=12'hA70;
20'b00000110010010011001:ColourData=12'hA70;
20'b00000110100010011001:ColourData=12'hC70;
20'b00000110110010011001:ColourData=12'hF93;
20'b00000111000010011001:ColourData=12'hF93;
20'b00000111010010011001:ColourData=12'hF93;
20'b00000111100010011001:ColourData=12'hAB2;
20'b00000111110010011001:ColourData=12'h8F7;
20'b00000000000010011010:ColourData=12'hC64;
20'b00000000010010011010:ColourData=12'hD72;
20'b00000000100010011010:ColourData=12'hE93;
20'b00000000110010011010:ColourData=12'hE83;
20'b00000001000010011010:ColourData=12'hE83;
20'b00000001010010011010:ColourData=12'hE83;
20'b00000001100010011010:ColourData=12'hE93;
20'b00000001110010011010:ColourData=12'hD72;
20'b00000010000010011010:ColourData=12'h310;
20'b00000010010010011010:ColourData=12'h210;
20'b00000010100010011010:ColourData=12'hD83;
20'b00000010110010011010:ColourData=12'hF93;
20'b00000011000010011010:ColourData=12'hE83;
20'b00000011010010011010:ColourData=12'hF93;
20'b00000011100010011010:ColourData=12'hC72;
20'b00000011110010011010:ColourData=12'h342;
20'b00000100000010011010:ColourData=12'h4F2;
20'b00000100010010011010:ColourData=12'h6C1;
20'b00000100100010011010:ColourData=12'hE30;
20'b00000100110010011010:ColourData=12'hF20;
20'b00000101000010011010:ColourData=12'hE30;
20'b00000101010010011010:ColourData=12'hB60;
20'b00000101100010011010:ColourData=12'hB60;
20'b00000101110010011010:ColourData=12'hB70;
20'b00000110000010011010:ColourData=12'hB50;
20'b00000110010010011010:ColourData=12'hA70;
20'b00000110100010011010:ColourData=12'h9A1;
20'b00000110110010011010:ColourData=12'hCB3;
20'b00000111000010011010:ColourData=12'hCB3;
20'b00000111010010011010:ColourData=12'hCB3;
20'b00000111100010011010:ColourData=12'h8C2;
20'b00000111110010011010:ColourData=12'h8F7;
20'b00000000000010011011:ColourData=12'hC64;
20'b00000000010010011011:ColourData=12'hD72;
20'b00000000100010011011:ColourData=12'hF93;
20'b00000000110010011011:ColourData=12'hE83;
20'b00000001000010011011:ColourData=12'hE83;
20'b00000001010010011011:ColourData=12'hE93;
20'b00000001100010011011:ColourData=12'hE83;
20'b00000001110010011011:ColourData=12'hC51;
20'b00000010000010011011:ColourData=12'hA41;
20'b00000010010010011011:ColourData=12'hC72;
20'b00000010100010011011:ColourData=12'hE83;
20'b00000010110010011011:ColourData=12'hE83;
20'b00000011000010011011:ColourData=12'hE83;
20'b00000011010010011011:ColourData=12'hF93;
20'b00000011100010011011:ColourData=12'hC72;
20'b00000011110010011011:ColourData=12'h342;
20'b00000100000010011011:ColourData=12'h4F2;
20'b00000100010010011011:ColourData=12'h6C1;
20'b00000100100010011011:ColourData=12'hE30;
20'b00000100110010011011:ColourData=12'hF20;
20'b00000101000010011011:ColourData=12'hF30;
20'b00000101010010011011:ColourData=12'hF20;
20'b00000101100010011011:ColourData=12'hF40;
20'b00000101110010011011:ColourData=12'hF61;
20'b00000110000010011011:ColourData=12'hF20;
20'b00000110010010011011:ColourData=12'hB60;
20'b00000110100010011011:ColourData=12'h3F1;
20'b00000110110010011011:ColourData=12'h3F1;
20'b00000111000010011011:ColourData=12'h4F1;
20'b00000111010010011011:ColourData=12'h5D1;
20'b00000111100010011011:ColourData=12'h4E0;
20'b00000111110010011011:ColourData=12'h8F7;
20'b00000000000010011100:ColourData=12'hC64;
20'b00000000010010011100:ColourData=12'hD72;
20'b00000000100010011100:ColourData=12'hD83;
20'b00000000110010011100:ColourData=12'hE83;
20'b00000001000010011100:ColourData=12'hE83;
20'b00000001010010011100:ColourData=12'hE93;
20'b00000001100010011100:ColourData=12'hE83;
20'b00000001110010011100:ColourData=12'hC51;
20'b00000010000010011100:ColourData=12'h931;
20'b00000010010010011100:ColourData=12'h310;
20'b00000010100010011100:ColourData=12'hD73;
20'b00000010110010011100:ColourData=12'hF93;
20'b00000011000010011100:ColourData=12'hE83;
20'b00000011010010011100:ColourData=12'hD83;
20'b00000011100010011100:ColourData=12'hC72;
20'b00000011110010011100:ColourData=12'h342;
20'b00000100000010011100:ColourData=12'h4F2;
20'b00000100010010011100:ColourData=12'h6C1;
20'b00000100100010011100:ColourData=12'hF20;
20'b00000100110010011100:ColourData=12'hF20;
20'b00000101000010011100:ColourData=12'hF30;
20'b00000101010010011100:ColourData=12'hF30;
20'b00000101100010011100:ColourData=12'hF30;
20'b00000101110010011100:ColourData=12'hF30;
20'b00000110000010011100:ColourData=12'hF20;
20'b00000110010010011100:ColourData=12'hC60;
20'b00000110100010011100:ColourData=12'h6C1;
20'b00000110110010011100:ColourData=12'h5C1;
20'b00000111000010011100:ColourData=12'h7B0;
20'b00000111010010011100:ColourData=12'hA60;
20'b00000111100010011100:ColourData=12'h7A0;
20'b00000111110010011100:ColourData=12'h8F7;
20'b00000000000010011101:ColourData=12'hC64;
20'b00000000010010011101:ColourData=12'hD72;
20'b00000000100010011101:ColourData=12'h531;
20'b00000000110010011101:ColourData=12'hC72;
20'b00000001000010011101:ColourData=12'hF93;
20'b00000001010010011101:ColourData=12'hE93;
20'b00000001100010011101:ColourData=12'hF93;
20'b00000001110010011101:ColourData=12'hE83;
20'b00000010000010011101:ColourData=12'h310;
20'b00000010010010011101:ColourData=12'h100;
20'b00000010100010011101:ColourData=12'hD83;
20'b00000010110010011101:ColourData=12'hF93;
20'b00000011000010011101:ColourData=12'hD83;
20'b00000011010010011101:ColourData=12'h531;
20'b00000011100010011101:ColourData=12'hB62;
20'b00000011110010011101:ColourData=12'h352;
20'b00000100000010011101:ColourData=12'h4F2;
20'b00000100010010011101:ColourData=12'h5D1;
20'b00000100100010011101:ColourData=12'hC50;
20'b00000100110010011101:ColourData=12'hF20;
20'b00000101000010011101:ColourData=12'hF30;
20'b00000101010010011101:ColourData=12'hF30;
20'b00000101100010011101:ColourData=12'hF30;
20'b00000101110010011101:ColourData=12'hF30;
20'b00000110000010011101:ColourData=12'hF30;
20'b00000110010010011101:ColourData=12'hE30;
20'b00000110100010011101:ColourData=12'hF30;
20'b00000110110010011101:ColourData=12'hD40;
20'b00000111000010011101:ColourData=12'hA70;
20'b00000111010010011101:ColourData=12'hA60;
20'b00000111100010011101:ColourData=12'h7A0;
20'b00000111110010011101:ColourData=12'h8F7;
20'b00000000000010011110:ColourData=12'hB64;
20'b00000000010010011110:ColourData=12'hC62;
20'b00000000100010011110:ColourData=12'hC72;
20'b00000000110010011110:ColourData=12'hC73;
20'b00000001000010011110:ColourData=12'hD83;
20'b00000001010010011110:ColourData=12'hD83;
20'b00000001100010011110:ColourData=12'hD83;
20'b00000001110010011110:ColourData=12'hD83;
20'b00000010000010011110:ColourData=12'hB72;
20'b00000010010010011110:ColourData=12'hB72;
20'b00000010100010011110:ColourData=12'hD73;
20'b00000010110010011110:ColourData=12'hD83;
20'b00000011000010011110:ColourData=12'hD73;
20'b00000011010010011110:ColourData=12'hC72;
20'b00000011100010011110:ColourData=12'hB62;
20'b00000011110010011110:ColourData=12'h342;
20'b00000100000010011110:ColourData=12'h4F1;
20'b00000100010010011110:ColourData=12'h3F1;
20'b00000100100010011110:ColourData=12'h5D0;
20'b00000100110010011110:ColourData=12'hC50;
20'b00000101000010011110:ColourData=12'hF20;
20'b00000101010010011110:ColourData=12'hF20;
20'b00000101100010011110:ColourData=12'hF20;
20'b00000101110010011110:ColourData=12'hF20;
20'b00000110000010011110:ColourData=12'hF20;
20'b00000110010010011110:ColourData=12'hF20;
20'b00000110100010011110:ColourData=12'hF20;
20'b00000110110010011110:ColourData=12'hD40;
20'b00000111000010011110:ColourData=12'hA70;
20'b00000111010010011110:ColourData=12'hA60;
20'b00000111100010011110:ColourData=12'h7A0;
20'b00000111110010011110:ColourData=12'h8F7;
20'b00000000000010011111:ColourData=12'h333;
20'b00000000010010011111:ColourData=12'h000;
20'b00000000100010011111:ColourData=12'h000;
20'b00000000110010011111:ColourData=12'h000;
20'b00000001000010011111:ColourData=12'h000;
20'b00000001010010011111:ColourData=12'h000;
20'b00000001100010011111:ColourData=12'h000;
20'b00000001110010011111:ColourData=12'h000;
20'b00000010000010011111:ColourData=12'h000;
20'b00000010010010011111:ColourData=12'h000;
20'b00000010100010011111:ColourData=12'h000;
20'b00000010110010011111:ColourData=12'h000;
20'b00000011000010011111:ColourData=12'h000;
20'b00000011010010011111:ColourData=12'h000;
20'b00000011100010011111:ColourData=12'h000;
20'b00000011110010011111:ColourData=12'h342;
20'b00000100000010011111:ColourData=12'h7F5;
20'b00000100010010011111:ColourData=12'h6F4;
20'b00000100100010011111:ColourData=12'h6F4;
20'b00000100110010011111:ColourData=12'h8D4;
20'b00000101000010011111:ColourData=12'hF53;
20'b00000101010010011111:ColourData=12'hF53;
20'b00000101100010011111:ColourData=12'hF53;
20'b00000101110010011111:ColourData=12'hF53;
20'b00000110000010011111:ColourData=12'hF53;
20'b00000110010010011111:ColourData=12'hF53;
20'b00000110100010011111:ColourData=12'hF53;
20'b00000110110010011111:ColourData=12'hD63;
20'b00000111000010011111:ColourData=12'hB93;
20'b00000111010010011111:ColourData=12'hB83;
20'b00000111100010011111:ColourData=12'h9B3;
20'b00000111110010011111:ColourData=12'hAF9;

default: ColourData = 12'h000;

endcase
end

endmodule