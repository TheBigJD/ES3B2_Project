module VGA_Draw(
    input Master_Clock_In, Reset_N_In,
    input Disp_Ena_In,
    input [9:0] Val_Col_In, Val_Row_In,
    input Up, Down,
    input Left, Right,
    
    output reg [3:0] Red = 4'h0, 
    output reg [3:0] Blue = 4'h0, 
    output reg [3:0] Green = 4'h0
);

parameter Pixels_Horiz = 640; //Num of Pixels in X axis
parameter Pixels_Vert  = 480; //Num of Pixels in Y axis

parameter EdgeWidth = 0;

reg [9:0] xPosition = 0; // Value is 1/2(Horiz Pixels + xWidth)
reg [9:0] yPosition = 0; // Value is 1/2(Vert Pixels + yWidth)

parameter yWidth = 30 ;// same as for xWidth 
parameter xWidth = 30 ;// random value i thought would be big enoguh to show up. if it's not increase it by a chunk

reg [3:0] Colour_Counter = 0;
reg [15:0] Clock_Div = 0;

//	reg [0:8] Pix_Red   [0:8][3:0];
//	reg [0:8] Pix_Blue  [0:8][3:0];
//	reg [0:8] Pix_Green [0:8][3:0];
//	reg [3:0] Red, Blue, Green;

wire [11:0] Colour_Data_Background;
wire [11:0] Colour_Data_Tank;

reg [9:0] Tank_XInput, Tank_YInput = 10'b0;	
reg [9:0] PrevX, PrevY = 10'b0;

reg [9:0] xDivPos, yDivPos;
reg [9:0] Tank_xDivPos, Tank_yDivPos, Tank_xDivPos_1, Tank_yDivPos_1;

reg [0:79] TankArray_1 = 80'b0;
reg [3:0] TankArray_X_1 = 4'b0;
reg TankArray_1_0, TankArray_1_1, TankArray_1_2, TankArray_1_3;

reg [0:79] TankArray_2 = 80'b0;
reg [3:0] TankArray_X_2 = 4'b0;
reg TankArray_2_0, TankArray_2_1, TankArray_2_2, TankArray_2_3;

reg [0:79] TankArray_3 = 80'b0;
reg [3:0] TankArray_X_3 = 4'b0;
reg TankArray_3_0, TankArray_3_1, TankArray_3_2, TankArray_3_3;

reg [0:79] TankArray_4 = 80'b0;
reg [3:0] TankArray_X_4 = 4'b0;
reg TankArray_4_0, TankArray_4_1, TankArray_4_2, TankArray_4_3;

//Bottle M4 (.Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Background));

TankImage M5 (.Master_Clock_In(Master_Clock_In), .xInput(Tank_XInput), .yInput(Tank_YInput), .ColourData(Colour_Data_Tank));

reg [0:79] MapArray [0:14];
reg [0:79] MapArrayData_Y = 80'b0;
reg [3:0]  MapArray_X = 4'b0;
reg MapArrayData_X_3, MapArrayData_X_2, MapArrayData_X_1, MapArrayData_X_0;



always @(posedge Master_Clock_In)	
	begin
		if (Reset_N_In == 0)
			begin
                Red   = 4'h0;     
                Blue  = 4'h0;
                Green = 4'h0;
    
                xPosition = 0;
                yPosition = 0;
            
			end
		else 
			begin
			// Need control for map choice here
                MapArray[ 0] = 80'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
                MapArray[ 1] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                MapArray[ 2] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                MapArray[ 3] = 80'b0000_0010_0010_0010_0010_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0010_0010_0010_0010_0000;
                MapArray[ 4] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                MapArray[ 5] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0010_0010_0010_0011_0010_0010_0011_0010_0011_0011_0000;
                MapArray[ 6] = 80'b0000_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0000;
                MapArray[ 7] = 80'b0000_0010_0010_0010_0010_0010_0011_0010_0010_0010_0010_0010_0010_0011_0010_0010_0010_0010_0010_0000;
                MapArray[ 8] = 80'b0000_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0000;
                MapArray[ 9] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0010_0010_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                MapArray[10] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                MapArray[11] = 80'b0000_0010_0010_0010_0010_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0010_0010_0010_0010_0000;
                MapArray[12] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                MapArray[13] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                MapArray[14] = 80'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

 
            if (Disp_Ena_In == 0)
                begin
                    Red 	= {4{1'b0}};
                    Blue 	= {4{1'b0}};
                    Green 	= {4{1'b0}};
                end
        
            else
                begin
                    if ((Val_Col_In <= Pixels_Vert) & (Val_Row_In <= Pixels_Horiz)) 
                        begin

////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                            //do not delete this. or i kill you.
                            // this is the bit that takes the x/y coordinates and shuffles them into the 20by15 array
                            // This will give the data for essentially 'What should we do with the tank at this point?
                            // We need to observe points at (x, y), (x+w, y), (x,y+w), (x+w, y+w) and make sure that these points
                            //      that the tank movement is limited if it reaches a point where the tank cant move through.
                            // This will allow the basis for the bullets too. If it hits a breakable block, we can change the reg's
                            //      value at this point to 4'h0, and the tank will behave differently than it would if it was 4'h2.
                            
                            xDivPos = ((Val_Row_In[9:5])%20);
                            yDivPos = ((Val_Col_In[9:5])%15);
                            
                            MapArrayData_Y   = MapArray[yDivPos];
                            MapArrayData_X_3 = MapArrayData_Y[4*xDivPos];
                            MapArrayData_X_2 = MapArrayData_Y[4*xDivPos + 1];
                            MapArrayData_X_1 = MapArrayData_Y[4*xDivPos + 2];
                            MapArrayData_X_0 = MapArrayData_Y[4*xDivPos + 3];
                            
                            MapArray_X = {MapArrayData_X_3, MapArrayData_X_2, MapArrayData_X_1, MapArrayData_X_0 };

                            if ((Val_Col_In == Pixels_Vert) & (Val_Row_In == Pixels_Horiz))
                                begin
////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                                    // If y-coordinate is at screen limit, move to other side of screen
                                    if (yPosition == EdgeWidth)
                                        yPosition = Pixels_Vert - yWidth;
                                    else if (yPosition == Pixels_Vert - yWidth - EdgeWidth)
                                        yPosition = 0;

                                    //if x-coordinate is at screen limit, move to other side of screen
                                    if (xPosition == EdgeWidth)
                                        xPosition = Pixels_Horiz - xWidth;
                                    else if (xPosition == Pixels_Horiz - xWidth - EdgeWidth)
                                        xPosition = 0;
////////////////////////////////////////////////////////////////////////////////////////////////////////////////                    
                                    //Setting Bounding boxes for tank control. Looking for box state at x and y positions
                                    Tank_xDivPos_1 = xPosition[9:5]%20;
                                    Tank_yDivPos_1 = yPosition[9:5]%15;
                                    
                                    Tank_xDivPos = ((xPosition + 20)/32)%20;
                                    Tank_yDivPos = ((yPosition + 20)/32)%15;
                                    
                                    
                                    //Bottom left
                                    TankArray_1   = MapArray[Tank_yDivPos_1];
                                    TankArray_1_3 = TankArray_1[4*Tank_xDivPos_1];
                                    TankArray_1_2 = TankArray_1[4*Tank_xDivPos_1+1];
                                    TankArray_1_1 = TankArray_1[4*Tank_xDivPos_1+2];
                                    TankArray_1_0 = TankArray_1[4*Tank_xDivPos_1+3];
                                    TankArray_X_1 = {TankArray_1_3,
 TankArray_1_2, TankArray_1_1, TankArray_1_0};
                                    //Bottom right
                                    TankArray_2   = MapArray[Tank_yDivPos_1];
                                    TankArray_2_3 = TankArray_2[4*(Tank_xDivPos )];
                                    TankArray_2_2 = TankArray_2[4*(Tank_xDivPos )+1];
                                    TankArray_2_1 = TankArray_2[4*(Tank_xDivPos )+2];
                                    TankArray_2_0 = TankArray_2[4*(Tank_xDivPos )+3];
                                    TankArray_X_2 = {TankArray_2_3, TankArray_2_2, TankArray_2_1, TankArray_2_0};   
                                    //Top left
                                    TankArray_3   = MapArray[Tank_yDivPos ];
                                    TankArray_3_3 = TankArray_3[4*(Tank_xDivPos_1)];
                                    TankArray_3_2 = TankArray_3[4*(Tank_xDivPos_1)+1];
                                    TankArray_3_1 = TankArray_3[4*(Tank_xDivPos_1)+2];
                                    TankArray_3_0 = TankArray_3[4*(Tank_xDivPos_1)+3];
                                    TankArray_X_3 = {TankArray_3_3, TankArray_3_2, TankArray_3_1, TankArray_3_0};   
                                    //Top right
                                    TankArray_4   = MapArray[Tank_yDivPos ];
                                    TankArray_4_3 = TankArray_4[4*(Tank_xDivPos)];
                                    TankArray_4_2 = TankArray_4[4*(Tank_xDivPos )+1];
                                    TankArray_4_1 = TankArray_4[4*(Tank_xDivPos )+2];
                                    TankArray_4_0 = TankArray_4[4*(Tank_xDivPos )+3];
                                    TankArray_X_4 = {TankArray_4_3, TankArray_4_2, TankArray_4_1, TankArray_4_0};                                    
                                    
                                    //If bottom edges are in boundary
                                            if ((TankArray_X_1 == 1) | (TankArray_X_1 == 2) | (TankArray_X_2 == 1) | (TankArray_X_2 == 2))
                                                yPosition = yPosition - 1;
                                    //If left edges are in boundary
                                    else    if ((TankArray_X_1 == 1) | (TankArray_X_1 == 2) | (TankArray_X_3 == 1) | (TankArray_X_3 == 2))
                                                xPosition = xPosition + 1;
                                    //if top edges are in boundary
                                    else    if ((TankArray_X_3 == 1) | (TankArray_X_3 == 2) | (TankArray_X_4 == 1) | (TankArray_X_4 == 2))
                                                yPosition = yPosition + 1;
                                    // if right edges are in boundary
                                    else    if ((TankArray_X_2 == 1) | (TankArray_X_2 == 2) | (TankArray_X_4 == 1) | (TankArray_X_4 == 2))
                                                xPosition = xPosition - 1;                        
                                 
                                end                                    
                                    
//                                    if ((TankArray_X_2 == 1) | (TankArray_X_2 == 2))
//                                        begin
//                                            yPosition = yPosition + 1;
//                                            xPosition = xPosition - 1;
//                                        end
//                                    else
//                                        begin
//                                            if (Up == 1)
//                                                yPosition = yPosition - 1;
//                                            if (Right == 1)
//                                                xPosition = xPosition + 1;

//                                            if ((TankArray_X_1 == 1) | (TankArray_X_1 == 2))
//                                                begin
//                                                    yPosition = yPosition - 1;
//                                                    xPosition = xPosition + 1;
//                                                end
//                                            else
//                                                begin
//                                                    if (Down == 1)
//                                                        yPosition = yPosition + 1;
//                                                    if (Left == 1)
//                                                        xPosition = xPosition - 1;
                                                        
//                                                end
//                                        end
//                                end     
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                            
                            
                            //within tank bounding box, set image to tank
                            if ((Val_Col_In >= yPosition) & (Val_Col_In <= yPosition + yWidth) & (Val_Row_In >= xPosition) & (Val_Row_In <= xPosition + xWidth))
                                begin
                                    PrevY = yPosition;
                                    PrevX = xPosition;
            
                                if (Down == 1)    
                                    begin
                                        Tank_XInput = xWidth - (Val_Row_In - xPosition)%xWidth;
                                        Tank_YInput = yWidth - (Val_Col_In - yPosition)%yWidth;
                                    end
            
                                else if (Left == 1)    
                                    begin
                                        Tank_YInput = Val_Row_In - xPosition;
                                        Tank_XInput = Val_Col_In - yPosition;
                                    end
            
                                else if (Right == 1)
                                    begin
                                        Tank_YInput = xWidth - (Val_Row_In - xPosition)%xWidth;
                                        Tank_XInput = yWidth - (Val_Col_In - yPosition)%yWidth;
                                    end
            
                                else
                                    begin
                                        Tank_XInput = Val_Row_In - xPosition;
                                        Tank_YInput = Val_Col_In - yPosition;
                                    end
            
            
                                    Red   = Colour_Data_Tank[11:8];
                                    Green = Colour_Data_Tank[7:4];
                                    Blue  = Colour_Data_Tank[3:0];
                                
                                end
                            else
                                //if not within tank bounding box
                                begin
            
    //                                if ((Val_Row_In <= EdgeWidth) | (Val_Row_In >= Pixels_Horiz - EdgeWidth) | (Val_Col_In <= EdgeWidth) | (Val_Col_In >= Pixels_Vert - EdgeWidth))
    //                                    begin
    //                                        Red 	= 4'h2;
    //                                        Green 	= 4'h2;
    //                                        Blue 	= 4'h2;
                                            
                                            
                                               
    ////                                        Red    = 4'h0;
    ////                                        Green  = 4'hF;
    ////                                        Blue   = 4'h0;
    //                                    end
    //                                else
                                       // begin
                                            
                                            //xDivPos = Val_Row_In[9:5]/32;
                                            //yDivPos = Val_Col_In[9:5]/32;
                                            
    
                                            case (MapArray_X)
                                                4'h0:begin  Red = 4'h0; Green = 4'h0; Blue = 4'hF; end
                                                4'h1:begin  Red = 4'h4; Green = 4'h4; Blue = 4'h4; end
                                                4'h2:begin  Red = 4'hF; Green = 4'h0; Blue = 4'h0; end
                                                4'h3:begin  Red = 4'hF; Green = 4'hF; Blue = 4'h0; end 
                                                
                                                default:begin Red = 4'h8; Green = 4'h8; Blue = 4'h8;end
                                                
                                            endcase
    //                                    end
            
                                end            
                    end
                
                else
                    begin
                        Red 	= 4'h2;
                        Blue 	= 4'h2;
                        Green 	= 4'h2;
                    end
                end
            end
        end

endmodule
