module MysteryImage(

  input Master_Clock_In,
  input [9 : 0] xInput,
  input [9 : 0] yInput,
  output reg [11:0] ColourData = 12'h000

);

(* rom_style = "block" *)

reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

always @(posedge Master_Clock_In)
begin
  a = xInput % 32;
  b = yInput % 32;

Inputs = {a, b};

    case(Inputs)
    //Converted_Image
20'b00000000000000000000 : ColourData = 12'hFFF;
20'b00000000010000000000 : ColourData = 12'hFFF;
20'b00000000100000000000 : ColourData = 12'hFFF;
20'b00000000110000000000 : ColourData = 12'hFFF;
20'b00000001000000000000 : ColourData = 12'hFFF;
20'b00000001010000000000 : ColourData = 12'hFFF;
20'b00000001100000000000 : ColourData = 12'hFFF;
20'b00000001110000000000 : ColourData = 12'hFFF;
20'b00000010000000000000 : ColourData = 12'hFFF;
20'b00000010010000000000 : ColourData = 12'hFFF;
20'b00000010100000000000 : ColourData = 12'hFFF;
20'b00000010110000000000 : ColourData = 12'hFFF;
20'b00000011000000000000 : ColourData = 12'hFFF;
20'b00000011010000000000 : ColourData = 12'hFFF;
20'b00000011100000000000 : ColourData = 12'hFFF;
20'b00000011110000000000 : ColourData = 12'hFFF;
20'b00000100000000000000 : ColourData = 12'hFFF;
20'b00000100010000000000 : ColourData = 12'hFFF;
20'b00000100100000000000 : ColourData = 12'hFFF;
20'b00000100110000000000 : ColourData = 12'hFFF;
20'b00000101000000000000 : ColourData = 12'hFFF;
20'b00000101010000000000 : ColourData = 12'hFFF;
20'b00000101100000000000 : ColourData = 12'hFFF;
20'b00000101110000000000 : ColourData = 12'hFFF;
20'b00000110000000000000 : ColourData = 12'hFFF;
20'b00000110010000000000 : ColourData = 12'hFFF;
20'b00000110100000000000 : ColourData = 12'hFFF;
20'b00000110110000000000 : ColourData = 12'hFFF;
20'b00000111000000000000 : ColourData = 12'hFFF;
20'b00000111010000000000 : ColourData = 12'hFFF;
20'b00000111100000000000 : ColourData = 12'hFFF;
20'b00000111110000000000 : ColourData = 12'hFFF;
20'b00000000000000000001 : ColourData = 12'hFFF;
20'b00000000010000000001 : ColourData = 12'hFFF;
20'b00000000100000000001 : ColourData = 12'hFFF;
20'b00000000110000000001 : ColourData = 12'hFFF;
20'b00000001000000000001 : ColourData = 12'hFFF;
20'b00000001010000000001 : ColourData = 12'hFFF;
20'b00000001100000000001 : ColourData = 12'hFFF;
20'b00000001110000000001 : ColourData = 12'hFFF;
20'b00000010000000000001 : ColourData = 12'hFFF;
20'b00000010010000000001 : ColourData = 12'hFFF;
20'b00000010100000000001 : ColourData = 12'hFFF;
20'b00000010110000000001 : ColourData = 12'hFFF;
20'b00000011000000000001 : ColourData = 12'hFFF;
20'b00000011010000000001 : ColourData = 12'hFFF;
20'b00000011100000000001 : ColourData = 12'hFFF;
20'b00000011110000000001 : ColourData = 12'hFFF;
20'b00000100000000000001 : ColourData = 12'hFFF;
20'b00000100010000000001 : ColourData = 12'hFFF;
20'b00000100100000000001 : ColourData = 12'hFFF;
20'b00000100110000000001 : ColourData = 12'hFFF;
20'b00000101000000000001 : ColourData = 12'hFFF;
20'b00000101010000000001 : ColourData = 12'hFFF;
20'b00000101100000000001 : ColourData = 12'hFFF;
20'b00000101110000000001 : ColourData = 12'hFFF;
20'b00000110000000000001 : ColourData = 12'hFFF;
20'b00000110010000000001 : ColourData = 12'hFFF;
20'b00000110100000000001 : ColourData = 12'hFFF;
20'b00000110110000000001 : ColourData = 12'hFFF;
20'b00000111000000000001 : ColourData = 12'hFFF;
20'b00000111010000000001 : ColourData = 12'hFFF;
20'b00000111100000000001 : ColourData = 12'hFFF;
20'b00000111110000000001 : ColourData = 12'hFFF;
20'b00000000000000000010 : ColourData = 12'hFFF;
20'b00000000010000000010 : ColourData = 12'hFFF;
20'b00000000100000000010 : ColourData = 12'hFFF;
20'b00000000110000000010 : ColourData = 12'hFFF;
20'b00000001000000000010 : ColourData = 12'hFFF;
20'b00000001010000000010 : ColourData = 12'hFFF;
20'b00000001100000000010 : ColourData = 12'hFFF;
20'b00000001110000000010 : ColourData = 12'hFFF;
20'b00000010000000000010 : ColourData = 12'hABB;
20'b00000010010000000010 : ColourData = 12'h9AA;
20'b00000010100000000010 : ColourData = 12'hAAA;
20'b00000010110000000010 : ColourData = 12'hAAA;
20'b00000011000000000010 : ColourData = 12'hAAA;
20'b00000011010000000010 : ColourData = 12'hAAA;
20'b00000011100000000010 : ColourData = 12'hAAA;
20'b00000011110000000010 : ColourData = 12'hAAA;
20'b00000100000000000010 : ColourData = 12'hAAB;
20'b00000100010000000010 : ColourData = 12'hAAB;
20'b00000100100000000010 : ColourData = 12'hBBB;
20'b00000100110000000010 : ColourData = 12'hBBB;
20'b00000101000000000010 : ColourData = 12'hBBB;
20'b00000101010000000010 : ColourData = 12'hBBB;
20'b00000101100000000010 : ColourData = 12'hBBB;
20'b00000101110000000010 : ColourData = 12'hBBC;
20'b00000110000000000010 : ColourData = 12'hFFF;
20'b00000110010000000010 : ColourData = 12'hFFF;
20'b00000110100000000010 : ColourData = 12'hFFF;
20'b00000110110000000010 : ColourData = 12'hFFF;
20'b00000111000000000010 : ColourData = 12'hFFF;
20'b00000111010000000010 : ColourData = 12'hFFF;
20'b00000111100000000010 : ColourData = 12'hFFF;
20'b00000111110000000010 : ColourData = 12'hFFF;
20'b00000000000000000011 : ColourData = 12'hFFF;
20'b00000000010000000011 : ColourData = 12'hFFF;
20'b00000000100000000011 : ColourData = 12'hFFF;
20'b00000000110000000011 : ColourData = 12'hFFF;
20'b00000001000000000011 : ColourData = 12'hFFF;
20'b00000001010000000011 : ColourData = 12'hFFF;
20'b00000001100000000011 : ColourData = 12'hFFF;
20'b00000001110000000011 : ColourData = 12'hFFF;
20'b00000010000000000011 : ColourData = 12'h222;
20'b00000010010000000011 : ColourData = 12'h000;
20'b00000010100000000011 : ColourData = 12'h000;
20'b00000010110000000011 : ColourData = 12'h000;
20'b00000011000000000011 : ColourData = 12'h000;
20'b00000011010000000011 : ColourData = 12'h000;
20'b00000011100000000011 : ColourData = 12'h000;
20'b00000011110000000011 : ColourData = 12'h000;
20'b00000100000000000011 : ColourData = 12'h000;
20'b00000100010000000011 : ColourData = 12'h000;
20'b00000100100000000011 : ColourData = 12'h000;
20'b00000100110000000011 : ColourData = 12'h000;
20'b00000101000000000011 : ColourData = 12'h000;
20'b00000101010000000011 : ColourData = 12'h000;
20'b00000101100000000011 : ColourData = 12'h000;
20'b00000101110000000011 : ColourData = 12'h001;
20'b00000110000000000011 : ColourData = 12'hEEE;
20'b00000110010000000011 : ColourData = 12'hFFF;
20'b00000110100000000011 : ColourData = 12'hFFF;
20'b00000110110000000011 : ColourData = 12'hFFF;
20'b00000111000000000011 : ColourData = 12'hFFF;
20'b00000111010000000011 : ColourData = 12'hFFF;
20'b00000111100000000011 : ColourData = 12'hFFF;
20'b00000111110000000011 : ColourData = 12'hFFF;
20'b00000000000000000100 : ColourData = 12'hFFF;
20'b00000000010000000100 : ColourData = 12'hFFF;
20'b00000000100000000100 : ColourData = 12'hFFF;
20'b00000000110000000100 : ColourData = 12'hFFF;
20'b00000001000000000100 : ColourData = 12'hFFF;
20'b00000001010000000100 : ColourData = 12'hFFF;
20'b00000001100000000100 : ColourData = 12'hFFF;
20'b00000001110000000100 : ColourData = 12'h999;
20'b00000010000000000100 : ColourData = 12'h985;
20'b00000010010000000100 : ColourData = 12'hB96;
20'b00000010100000000100 : ColourData = 12'hB96;
20'b00000010110000000100 : ColourData = 12'hB96;
20'b00000011000000000100 : ColourData = 12'hB96;
20'b00000011010000000100 : ColourData = 12'hB96;
20'b00000011100000000100 : ColourData = 12'hB96;
20'b00000011110000000100 : ColourData = 12'hB96;
20'b00000100000000000100 : ColourData = 12'hB96;
20'b00000100010000000100 : ColourData = 12'hB96;
20'b00000100100000000100 : ColourData = 12'hB96;
20'b00000100110000000100 : ColourData = 12'hB96;
20'b00000101000000000100 : ColourData = 12'hB96;
20'b00000101010000000100 : ColourData = 12'hB96;
20'b00000101100000000100 : ColourData = 12'hB96;
20'b00000101110000000100 : ColourData = 12'hA86;
20'b00000110000000000100 : ColourData = 12'h666;
20'b00000110010000000100 : ColourData = 12'hFFF;
20'b00000110100000000100 : ColourData = 12'hFFF;
20'b00000110110000000100 : ColourData = 12'hFFF;
20'b00000111000000000100 : ColourData = 12'hFFF;
20'b00000111010000000100 : ColourData = 12'hFFF;
20'b00000111100000000100 : ColourData = 12'hFFF;
20'b00000111110000000100 : ColourData = 12'hFFF;
20'b00000000000000000101 : ColourData = 12'hFFF;
20'b00000000010000000101 : ColourData = 12'hFFF;
20'b00000000100000000101 : ColourData = 12'hFFF;
20'b00000000110000000101 : ColourData = 12'hFFF;
20'b00000001000000000101 : ColourData = 12'hFFF;
20'b00000001010000000101 : ColourData = 12'hFFF;
20'b00000001100000000101 : ColourData = 12'h999;
20'b00000001110000000101 : ColourData = 12'h765;
20'b00000010000000000101 : ColourData = 12'hEB8;
20'b00000010010000000101 : ColourData = 12'hFC9;
20'b00000010100000000101 : ColourData = 12'hFAC;
20'b00000010110000000101 : ColourData = 12'hFAD;
20'b00000011000000000101 : ColourData = 12'hFAD;
20'b00000011010000000101 : ColourData = 12'hFAD;
20'b00000011100000000101 : ColourData = 12'hFAD;
20'b00000011110000000101 : ColourData = 12'hFAD;
20'b00000100000000000101 : ColourData = 12'hFAD;
20'b00000100010000000101 : ColourData = 12'hFAD;
20'b00000100100000000101 : ColourData = 12'hFAD;
20'b00000100110000000101 : ColourData = 12'hFAD;
20'b00000101000000000101 : ColourData = 12'hFAD;
20'b00000101010000000101 : ColourData = 12'hFAC;
20'b00000101100000000101 : ColourData = 12'hFC9;
20'b00000101110000000101 : ColourData = 12'hFC8;
20'b00000110000000000101 : ColourData = 12'h875;
20'b00000110010000000101 : ColourData = 12'h889;
20'b00000110100000000101 : ColourData = 12'hFFF;
20'b00000110110000000101 : ColourData = 12'hFFF;
20'b00000111000000000101 : ColourData = 12'hFFF;
20'b00000111010000000101 : ColourData = 12'hFFF;
20'b00000111100000000101 : ColourData = 12'hFFF;
20'b00000111110000000101 : ColourData = 12'hFFF;
20'b00000000000000000110 : ColourData = 12'hFFF;
20'b00000000010000000110 : ColourData = 12'hFFF;
20'b00000000100000000110 : ColourData = 12'hFFF;
20'b00000000110000000110 : ColourData = 12'hFFF;
20'b00000001000000000110 : ColourData = 12'hFFF;
20'b00000001010000000110 : ColourData = 12'hFFF;
20'b00000001100000000110 : ColourData = 12'h444;
20'b00000001110000000110 : ColourData = 12'h864;
20'b00000010000000000110 : ColourData = 12'hFD9;
20'b00000010010000000110 : ColourData = 12'hFB9;
20'b00000010100000000110 : ColourData = 12'hF9E;
20'b00000010110000000110 : ColourData = 12'hF8F;
20'b00000011000000000110 : ColourData = 12'hF8F;
20'b00000011010000000110 : ColourData = 12'hF8F;
20'b00000011100000000110 : ColourData = 12'hF8F;
20'b00000011110000000110 : ColourData = 12'hF8F;
20'b00000100000000000110 : ColourData = 12'hF8F;
20'b00000100010000000110 : ColourData = 12'hF8F;
20'b00000100100000000110 : ColourData = 12'hF8F;
20'b00000100110000000110 : ColourData = 12'hF8F;
20'b00000101000000000110 : ColourData = 12'hF8F;
20'b00000101010000000110 : ColourData = 12'hF8F;
20'b00000101100000000110 : ColourData = 12'hFBA;
20'b00000101110000000110 : ColourData = 12'hFC9;
20'b00000110000000000110 : ColourData = 12'hCA7;
20'b00000110010000000110 : ColourData = 12'h333;
20'b00000110100000000110 : ColourData = 12'hFFF;
20'b00000110110000000110 : ColourData = 12'hFFF;
20'b00000111000000000110 : ColourData = 12'hFFF;
20'b00000111010000000110 : ColourData = 12'hFFF;
20'b00000111100000000110 : ColourData = 12'hFFF;
20'b00000111110000000110 : ColourData = 12'hFFF;
20'b00000000000000000111 : ColourData = 12'hFFF;
20'b00000000010000000111 : ColourData = 12'hFFF;
20'b00000000100000000111 : ColourData = 12'hFFF;
20'b00000000110000000111 : ColourData = 12'hFFF;
20'b00000001000000000111 : ColourData = 12'hFFF;
20'b00000001010000000111 : ColourData = 12'hFFF;
20'b00000001100000000111 : ColourData = 12'h455;
20'b00000001110000000111 : ColourData = 12'h864;
20'b00000010000000000111 : ColourData = 12'hFC9;
20'b00000010010000000111 : ColourData = 12'hF9D;
20'b00000010100000000111 : ColourData = 12'hF9F;
20'b00000010110000000111 : ColourData = 12'hF8F;
20'b00000011000000000111 : ColourData = 12'hF8F;
20'b00000011010000000111 : ColourData = 12'hF9F;
20'b00000011100000000111 : ColourData = 12'hF5C;
20'b00000011110000000111 : ColourData = 12'hF4B;
20'b00000100000000000111 : ColourData = 12'hF9F;
20'b00000100010000000111 : ColourData = 12'hF5C;
20'b00000100100000000111 : ColourData = 12'hF6C;
20'b00000100110000000111 : ColourData = 12'hF9F;
20'b00000101000000000111 : ColourData = 12'hF8F;
20'b00000101010000000111 : ColourData = 12'hF8F;
20'b00000101100000000111 : ColourData = 12'hF9E;
20'b00000101110000000111 : ColourData = 12'hFC9;
20'b00000110000000000111 : ColourData = 12'hCA7;
20'b00000110010000000111 : ColourData = 12'h444;
20'b00000110100000000111 : ColourData = 12'hFFF;
20'b00000110110000000111 : ColourData = 12'hFFF;
20'b00000111000000000111 : ColourData = 12'hFFF;
20'b00000111010000000111 : ColourData = 12'hFFF;
20'b00000111100000000111 : ColourData = 12'hFFF;
20'b00000111110000000111 : ColourData = 12'hFFF;
20'b00000000000000001000 : ColourData = 12'hFFF;
20'b00000000010000001000 : ColourData = 12'hFFF;
20'b00000000100000001000 : ColourData = 12'hFFF;
20'b00000000110000001000 : ColourData = 12'hEBB;
20'b00000001000000001000 : ColourData = 12'hE99;
20'b00000001010000001000 : ColourData = 12'hE99;
20'b00000001100000001000 : ColourData = 12'h423;
20'b00000001110000001000 : ColourData = 12'h874;
20'b00000010000000001000 : ColourData = 12'hFBB;
20'b00000010010000001000 : ColourData = 12'hF8E;
20'b00000010100000001000 : ColourData = 12'hF5C;
20'b00000010110000001000 : ColourData = 12'hF8E;
20'b00000011000000001000 : ColourData = 12'hF8F;
20'b00000011010000001000 : ColourData = 12'hF9F;
20'b00000011100000001000 : ColourData = 12'hF7D;
20'b00000011110000001000 : ColourData = 12'hF6D;
20'b00000100000000001000 : ColourData = 12'hF9F;
20'b00000100010000001000 : ColourData = 12'hF7E;
20'b00000100100000001000 : ColourData = 12'hF7E;
20'b00000100110000001000 : ColourData = 12'hF9F;
20'b00000101000000001000 : ColourData = 12'hF8F;
20'b00000101010000001000 : ColourData = 12'hF8F;
20'b00000101100000001000 : ColourData = 12'hF8F;
20'b00000101110000001000 : ColourData = 12'hFAC;
20'b00000110000000001000 : ColourData = 12'hC97;
20'b00000110010000001000 : ColourData = 12'h444;
20'b00000110100000001000 : ColourData = 12'hFFF;
20'b00000110110000001000 : ColourData = 12'hFFF;
20'b00000111000000001000 : ColourData = 12'hFFF;
20'b00000111010000001000 : ColourData = 12'hFFF;
20'b00000111100000001000 : ColourData = 12'hFFF;
20'b00000111110000001000 : ColourData = 12'hFFF;
20'b00000000000000001001 : ColourData = 12'hEFF;
20'b00000000010000001001 : ColourData = 12'hEFF;
20'b00000000100000001001 : ColourData = 12'hEFF;
20'b00000000110000001001 : ColourData = 12'hE23;
20'b00000001000000001001 : ColourData = 12'hF00;
20'b00000001010000001001 : ColourData = 12'hF00;
20'b00000001100000001001 : ColourData = 12'h400;
20'b00000001110000001001 : ColourData = 12'h875;
20'b00000010000000001001 : ColourData = 12'hF9E;
20'b00000010010000001001 : ColourData = 12'hF8F;
20'b00000010100000001001 : ColourData = 12'hE3A;
20'b00000010110000001001 : ColourData = 12'hF8E;
20'b00000011000000001001 : ColourData = 12'hF9F;
20'b00000011010000001001 : ColourData = 12'hF8F;
20'b00000011100000001001 : ColourData = 12'hF9F;
20'b00000011110000001001 : ColourData = 12'hF9F;
20'b00000100000000001001 : ColourData = 12'hF8F;
20'b00000100010000001001 : ColourData = 12'hE8E;
20'b00000100100000001001 : ColourData = 12'hE8E;
20'b00000100110000001001 : ColourData = 12'hF8F;
20'b00000101000000001001 : ColourData = 12'hF8F;
20'b00000101010000001001 : ColourData = 12'hF8E;
20'b00000101100000001001 : ColourData = 12'hF8F;
20'b00000101110000001001 : ColourData = 12'hF9F;
20'b00000110000000001001 : ColourData = 12'hC97;
20'b00000110010000001001 : ColourData = 12'h444;
20'b00000110100000001001 : ColourData = 12'hFFF;
20'b00000110110000001001 : ColourData = 12'hEEE;
20'b00000111000000001001 : ColourData = 12'hFFF;
20'b00000111010000001001 : ColourData = 12'hFFF;
20'b00000111100000001001 : ColourData = 12'hFFF;
20'b00000111110000001001 : ColourData = 12'hFFF;
20'b00000000000000001010 : ColourData = 12'hD22;
20'b00000000010000001010 : ColourData = 12'hD22;
20'b00000000100000001010 : ColourData = 12'hD22;
20'b00000000110000001010 : ColourData = 12'hE00;
20'b00000001000000001010 : ColourData = 12'hF00;
20'b00000001010000001010 : ColourData = 12'hF00;
20'b00000001100000001010 : ColourData = 12'h500;
20'b00000001110000001010 : ColourData = 12'h875;
20'b00000010000000001010 : ColourData = 12'hFAE;
20'b00000010010000001010 : ColourData = 12'hF8F;
20'b00000010100000001010 : ColourData = 12'hF8E;
20'b00000010110000001010 : ColourData = 12'hF8F;
20'b00000011000000001010 : ColourData = 12'hF8F;
20'b00000011010000001010 : ColourData = 12'hF8F;
20'b00000011100000001010 : ColourData = 12'hF8F;
20'b00000011110000001010 : ColourData = 12'hF8F;
20'b00000100000000001010 : ColourData = 12'hF9F;
20'b00000100010000001010 : ColourData = 12'h959;
20'b00000100100000001010 : ColourData = 12'h000;
20'b00000100110000001010 : ColourData = 12'hA6A;
20'b00000101000000001010 : ColourData = 12'hF9F;
20'b00000101010000001010 : ColourData = 12'hE3A;
20'b00000101100000001010 : ColourData = 12'hF7E;
20'b00000101110000001010 : ColourData = 12'hF9F;
20'b00000110000000001010 : ColourData = 12'hC97;
20'b00000110010000001010 : ColourData = 12'h444;
20'b00000110100000001010 : ColourData = 12'hEEE;
20'b00000110110000001010 : ColourData = 12'h222;
20'b00000111000000001010 : ColourData = 12'h666;
20'b00000111010000001010 : ColourData = 12'hFFF;
20'b00000111100000001010 : ColourData = 12'hFFF;
20'b00000111110000001010 : ColourData = 12'hFFF;
20'b00000000000000001011 : ColourData = 12'hF00;
20'b00000000010000001011 : ColourData = 12'hF00;
20'b00000000100000001011 : ColourData = 12'hF00;
20'b00000000110000001011 : ColourData = 12'hF10;
20'b00000001000000001011 : ColourData = 12'hF20;
20'b00000001010000001011 : ColourData = 12'hF20;
20'b00000001100000001011 : ColourData = 12'h500;
20'b00000001110000001011 : ColourData = 12'h875;
20'b00000010000000001011 : ColourData = 12'hFAE;
20'b00000010010000001011 : ColourData = 12'hF8F;
20'b00000010100000001011 : ColourData = 12'hF8F;
20'b00000010110000001011 : ColourData = 12'hF8F;
20'b00000011000000001011 : ColourData = 12'hF8F;
20'b00000011010000001011 : ColourData = 12'hF8F;
20'b00000011100000001011 : ColourData = 12'hF9F;
20'b00000011110000001011 : ColourData = 12'hF9F;
20'b00000100000000001011 : ColourData = 12'h959;
20'b00000100010000001011 : ColourData = 12'h434;
20'b00000100100000001011 : ColourData = 12'h777;
20'b00000100110000001011 : ColourData = 12'h333;
20'b00000101000000001011 : ColourData = 12'hA6A;
20'b00000101010000001011 : ColourData = 12'hF8E;
20'b00000101100000001011 : ColourData = 12'hF8F;
20'b00000101110000001011 : ColourData = 12'hF9F;
20'b00000110000000001011 : ColourData = 12'hCA7;
20'b00000110010000001011 : ColourData = 12'h000;
20'b00000110100000001011 : ColourData = 12'h333;
20'b00000110110000001011 : ColourData = 12'h777;
20'b00000111000000001011 : ColourData = 12'h555;
20'b00000111010000001011 : ColourData = 12'h999;
20'b00000111100000001011 : ColourData = 12'hFFF;
20'b00000111110000001011 : ColourData = 12'hFFF;
20'b00000000000000001100 : ColourData = 12'hE00;
20'b00000000010000001100 : ColourData = 12'hB00;
20'b00000000100000001100 : ColourData = 12'hA00;
20'b00000000110000001100 : ColourData = 12'hA50;
20'b00000001000000001100 : ColourData = 12'hC80;
20'b00000001010000001100 : ColourData = 12'hF90;
20'b00000001100000001100 : ColourData = 12'h520;
20'b00000001110000001100 : ColourData = 12'h875;
20'b00000010000000001100 : ColourData = 12'hFAE;
20'b00000010010000001100 : ColourData = 12'hF8F;
20'b00000010100000001100 : ColourData = 12'hF8F;
20'b00000010110000001100 : ColourData = 12'hF8F;
20'b00000011000000001100 : ColourData = 12'hF8F;
20'b00000011010000001100 : ColourData = 12'hF8E;
20'b00000011100000001100 : ColourData = 12'hF7E;
20'b00000011110000001100 : ColourData = 12'hF9F;
20'b00000100000000001100 : ColourData = 12'h848;
20'b00000100010000001100 : ColourData = 12'h232;
20'b00000100100000001100 : ColourData = 12'h999;
20'b00000100110000001100 : ColourData = 12'h444;
20'b00000101000000001100 : ColourData = 12'h747;
20'b00000101010000001100 : ColourData = 12'hE8E;
20'b00000101100000001100 : ColourData = 12'hF8F;
20'b00000101110000001100 : ColourData = 12'hF9F;
20'b00000110000000001100 : ColourData = 12'hCA8;
20'b00000110010000001100 : ColourData = 12'h000;
20'b00000110100000001100 : ColourData = 12'h222;
20'b00000110110000001100 : ColourData = 12'h999;
20'b00000111000000001100 : ColourData = 12'h555;
20'b00000111010000001100 : ColourData = 12'h777;
20'b00000111100000001100 : ColourData = 12'hFFF;
20'b00000111110000001100 : ColourData = 12'hFFF;
20'b00000000000000001101 : ColourData = 12'hC50;
20'b00000000010000001101 : ColourData = 12'h000;
20'b00000000100000001101 : ColourData = 12'h000;
20'b00000000110000001101 : ColourData = 12'h000;
20'b00000001000000001101 : ColourData = 12'h530;
20'b00000001010000001101 : ColourData = 12'hF90;
20'b00000001100000001101 : ColourData = 12'h520;
20'b00000001110000001101 : ColourData = 12'h875;
20'b00000010000000001101 : ColourData = 12'hFAE;
20'b00000010010000001101 : ColourData = 12'hF8F;
20'b00000010100000001101 : ColourData = 12'hF8F;
20'b00000010110000001101 : ColourData = 12'hF8F;
20'b00000011000000001101 : ColourData = 12'hF9F;
20'b00000011010000001101 : ColourData = 12'hF7D;
20'b00000011100000001101 : ColourData = 12'hF4B;
20'b00000011110000001101 : ColourData = 12'hF9F;
20'b00000100000000001101 : ColourData = 12'h848;
20'b00000100010000001101 : ColourData = 12'h333;
20'b00000100100000001101 : ColourData = 12'h999;
20'b00000100110000001101 : ColourData = 12'h999;
20'b00000101000000001101 : ColourData = 12'h333;
20'b00000101010000001101 : ColourData = 12'hC7C;
20'b00000101100000001101 : ColourData = 12'hF9F;
20'b00000101110000001101 : ColourData = 12'hF9F;
20'b00000110000000001101 : ColourData = 12'hCA8;
20'b00000110010000001101 : ColourData = 12'h222;
20'b00000110100000001101 : ColourData = 12'h999;
20'b00000110110000001101 : ColourData = 12'h999;
20'b00000111000000001101 : ColourData = 12'h555;
20'b00000111010000001101 : ColourData = 12'h777;
20'b00000111100000001101 : ColourData = 12'hFFF;
20'b00000111110000001101 : ColourData = 12'hFFF;
20'b00000000000000001110 : ColourData = 12'hC70;
20'b00000000010000001110 : ColourData = 12'h222;
20'b00000000100000001110 : ColourData = 12'h777;
20'b00000000110000001110 : ColourData = 12'h222;
20'b00000001000000001110 : ColourData = 12'h100;
20'b00000001010000001110 : ColourData = 12'hC80;
20'b00000001100000001110 : ColourData = 12'h530;
20'b00000001110000001110 : ColourData = 12'h875;
20'b00000010000000001110 : ColourData = 12'hFAE;
20'b00000010010000001110 : ColourData = 12'hF8F;
20'b00000010100000001110 : ColourData = 12'hF8F;
20'b00000010110000001110 : ColourData = 12'hF9F;
20'b00000011000000001110 : ColourData = 12'hF8F;
20'b00000011010000001110 : ColourData = 12'hF8E;
20'b00000011100000001110 : ColourData = 12'hF7E;
20'b00000011110000001110 : ColourData = 12'hF9F;
20'b00000100000000001110 : ColourData = 12'h848;
20'b00000100010000001110 : ColourData = 12'h333;
20'b00000100100000001110 : ColourData = 12'h999;
20'b00000100110000001110 : ColourData = 12'h999;
20'b00000101000000001110 : ColourData = 12'h777;
20'b00000101010000001110 : ColourData = 12'h424;
20'b00000101100000001110 : ColourData = 12'h323;
20'b00000101110000001110 : ColourData = 12'h323;
20'b00000110000000001110 : ColourData = 12'h432;
20'b00000110010000001110 : ColourData = 12'h777;
20'b00000110100000001110 : ColourData = 12'h999;
20'b00000110110000001110 : ColourData = 12'h999;
20'b00000111000000001110 : ColourData = 12'h555;
20'b00000111010000001110 : ColourData = 12'h777;
20'b00000111100000001110 : ColourData = 12'hFFF;
20'b00000111110000001110 : ColourData = 12'hFFF;
20'b00000000000000001111 : ColourData = 12'hC70;
20'b00000000010000001111 : ColourData = 12'h111;
20'b00000000100000001111 : ColourData = 12'h666;
20'b00000000110000001111 : ColourData = 12'h777;
20'b00000001000000001111 : ColourData = 12'h222;
20'b00000001010000001111 : ColourData = 12'h330;
20'b00000001100000001111 : ColourData = 12'h220;
20'b00000001110000001111 : ColourData = 12'h875;
20'b00000010000000001111 : ColourData = 12'hFAE;
20'b00000010010000001111 : ColourData = 12'hF8F;
20'b00000010100000001111 : ColourData = 12'hF8F;
20'b00000010110000001111 : ColourData = 12'hF5C;
20'b00000011000000001111 : ColourData = 12'hF8F;
20'b00000011010000001111 : ColourData = 12'hF8F;
20'b00000011100000001111 : ColourData = 12'hF9F;
20'b00000011110000001111 : ColourData = 12'hF9F;
20'b00000100000000001111 : ColourData = 12'h848;
20'b00000100010000001111 : ColourData = 12'h232;
20'b00000100100000001111 : ColourData = 12'h999;
20'b00000100110000001111 : ColourData = 12'h999;
20'b00000101000000001111 : ColourData = 12'h999;
20'b00000101010000001111 : ColourData = 12'h555;
20'b00000101100000001111 : ColourData = 12'h444;
20'b00000101110000001111 : ColourData = 12'h444;
20'b00000110000000001111 : ColourData = 12'h555;
20'b00000110010000001111 : ColourData = 12'h999;
20'b00000110100000001111 : ColourData = 12'h999;
20'b00000110110000001111 : ColourData = 12'h999;
20'b00000111000000001111 : ColourData = 12'h555;
20'b00000111010000001111 : ColourData = 12'h777;
20'b00000111100000001111 : ColourData = 12'hFFF;
20'b00000111110000001111 : ColourData = 12'hFFF;
20'b00000000000000010000 : ColourData = 12'hCA0;
20'b00000000010000010000 : ColourData = 12'h000;
20'b00000000100000010000 : ColourData = 12'h222;
20'b00000000110000010000 : ColourData = 12'h999;
20'b00000001000000010000 : ColourData = 12'h666;
20'b00000001010000010000 : ColourData = 12'h000;
20'b00000001100000010000 : ColourData = 12'h000;
20'b00000001110000010000 : ColourData = 12'h975;
20'b00000010000000010000 : ColourData = 12'hFAE;
20'b00000010010000010000 : ColourData = 12'hF8F;
20'b00000010100000010000 : ColourData = 12'hF8E;
20'b00000010110000010000 : ColourData = 12'hF3A;
20'b00000011000000010000 : ColourData = 12'hF8F;
20'b00000011010000010000 : ColourData = 12'hF8F;
20'b00000011100000010000 : ColourData = 12'hF8F;
20'b00000011110000010000 : ColourData = 12'hE8E;
20'b00000100000000010000 : ColourData = 12'h748;
20'b00000100010000010000 : ColourData = 12'h333;
20'b00000100100000010000 : ColourData = 12'h999;
20'b00000100110000010000 : ColourData = 12'h999;
20'b00000101000000010000 : ColourData = 12'h999;
20'b00000101010000010000 : ColourData = 12'h999;
20'b00000101100000010000 : ColourData = 12'h999;
20'b00000101110000010000 : ColourData = 12'h999;
20'b00000110000000010000 : ColourData = 12'h999;
20'b00000110010000010000 : ColourData = 12'h999;
20'b00000110100000010000 : ColourData = 12'h999;
20'b00000110110000010000 : ColourData = 12'h999;
20'b00000111000000010000 : ColourData = 12'h555;
20'b00000111010000010000 : ColourData = 12'h666;
20'b00000111100000010000 : ColourData = 12'hEEF;
20'b00000111110000010000 : ColourData = 12'hFFF;
20'b00000000000000010001 : ColourData = 12'hFF0;
20'b00000000010000010001 : ColourData = 12'h770;
20'b00000000100000010001 : ColourData = 12'h000;
20'b00000000110000010001 : ColourData = 12'h555;
20'b00000001000000010001 : ColourData = 12'h999;
20'b00000001010000010001 : ColourData = 12'h222;
20'b00000001100000010001 : ColourData = 12'h000;
20'b00000001110000010001 : ColourData = 12'h975;
20'b00000010000000010001 : ColourData = 12'hFAE;
20'b00000010010000010001 : ColourData = 12'hF8F;
20'b00000010100000010001 : ColourData = 12'hF8F;
20'b00000010110000010001 : ColourData = 12'hF8E;
20'b00000011000000010001 : ColourData = 12'hF8F;
20'b00000011010000010001 : ColourData = 12'hF9F;
20'b00000011100000010001 : ColourData = 12'hF6D;
20'b00000011110000010001 : ColourData = 12'h815;
20'b00000100000000010001 : ColourData = 12'h333;
20'b00000100010000010001 : ColourData = 12'h898;
20'b00000100100000010001 : ColourData = 12'h999;
20'b00000100110000010001 : ColourData = 12'h888;
20'b00000101000000010001 : ColourData = 12'h999;
20'b00000101010000010001 : ColourData = 12'h999;
20'b00000101100000010001 : ColourData = 12'h999;
20'b00000101110000010001 : ColourData = 12'h999;
20'b00000110000000010001 : ColourData = 12'h999;
20'b00000110010000010001 : ColourData = 12'h999;
20'b00000110100000010001 : ColourData = 12'h888;
20'b00000110110000010001 : ColourData = 12'h999;
20'b00000111000000010001 : ColourData = 12'h999;
20'b00000111010000010001 : ColourData = 12'h444;
20'b00000111100000010001 : ColourData = 12'h788;
20'b00000111110000010001 : ColourData = 12'hFFF;
20'b00000000000000010010 : ColourData = 12'hFF0;
20'b00000000010000010010 : ColourData = 12'hDD0;
20'b00000000100000010010 : ColourData = 12'h550;
20'b00000000110000010010 : ColourData = 12'h111;
20'b00000001000000010010 : ColourData = 12'h555;
20'b00000001010000010010 : ColourData = 12'h777;
20'b00000001100000010010 : ColourData = 12'h111;
20'b00000001110000010010 : ColourData = 12'h875;
20'b00000010000000010010 : ColourData = 12'hF9E;
20'b00000010010000010010 : ColourData = 12'hF5C;
20'b00000010100000010010 : ColourData = 12'hF8E;
20'b00000010110000010010 : ColourData = 12'hF9F;
20'b00000011000000010010 : ColourData = 12'hF8F;
20'b00000011010000010010 : ColourData = 12'hF8F;
20'b00000011100000010010 : ColourData = 12'hF8E;
20'b00000011110000010010 : ColourData = 12'h836;
20'b00000100000000010010 : ColourData = 12'h333;
20'b00000100010000010010 : ColourData = 12'h999;
20'b00000100100000010010 : ColourData = 12'h888;
20'b00000100110000010010 : ColourData = 12'hBBB;
20'b00000101000000010010 : ColourData = 12'h777;
20'b00000101010000010010 : ColourData = 12'h777;
20'b00000101100000010010 : ColourData = 12'h999;
20'b00000101110000010010 : ColourData = 12'h999;
20'b00000110000000010010 : ColourData = 12'h999;
20'b00000110010000010010 : ColourData = 12'hAAA;
20'b00000110100000010010 : ColourData = 12'hBBB;
20'b00000110110000010010 : ColourData = 12'h666;
20'b00000111000000010010 : ColourData = 12'h999;
20'b00000111010000010010 : ColourData = 12'h444;
20'b00000111100000010010 : ColourData = 12'h667;
20'b00000111110000010010 : ColourData = 12'hFFF;
20'b00000000000000010011 : ColourData = 12'h8F0;
20'b00000000010000010011 : ColourData = 12'h8F0;
20'b00000000100000010011 : ColourData = 12'h590;
20'b00000000110000010011 : ColourData = 12'h000;
20'b00000001000000010011 : ColourData = 12'h333;
20'b00000001010000010011 : ColourData = 12'h999;
20'b00000001100000010011 : ColourData = 12'h223;
20'b00000001110000010011 : ColourData = 12'h875;
20'b00000010000000010011 : ColourData = 12'hF9E;
20'b00000010010000010011 : ColourData = 12'hE3A;
20'b00000010100000010011 : ColourData = 12'hF8E;
20'b00000010110000010011 : ColourData = 12'hF9F;
20'b00000011000000010011 : ColourData = 12'hF8F;
20'b00000011010000010011 : ColourData = 12'hF8F;
20'b00000011100000010011 : ColourData = 12'hF9F;
20'b00000011110000010011 : ColourData = 12'h848;
20'b00000100000000010011 : ColourData = 12'h333;
20'b00000100010000010011 : ColourData = 12'h999;
20'b00000100100000010011 : ColourData = 12'h888;
20'b00000100110000010011 : ColourData = 12'hDDD;
20'b00000101000000010011 : ColourData = 12'h555;
20'b00000101010000010011 : ColourData = 12'h777;
20'b00000101100000010011 : ColourData = 12'h999;
20'b00000101110000010011 : ColourData = 12'h999;
20'b00000110000000010011 : ColourData = 12'h888;
20'b00000110010000010011 : ColourData = 12'hAAA;
20'b00000110100000010011 : ColourData = 12'hCCC;
20'b00000110110000010011 : ColourData = 12'h444;
20'b00000111000000010011 : ColourData = 12'h999;
20'b00000111010000010011 : ColourData = 12'h444;
20'b00000111100000010011 : ColourData = 12'h777;
20'b00000111110000010011 : ColourData = 12'hFFF;
20'b00000000000000010100 : ColourData = 12'h0F0;
20'b00000000010000010100 : ColourData = 12'h0F0;
20'b00000000100000010100 : ColourData = 12'h0E0;
20'b00000000110000010100 : ColourData = 12'h060;
20'b00000001000000010100 : ColourData = 12'h000;
20'b00000001010000010100 : ColourData = 12'h111;
20'b00000001100000010100 : ColourData = 12'h000;
20'b00000001110000010100 : ColourData = 12'h875;
20'b00000010000000010100 : ColourData = 12'hFAE;
20'b00000010010000010100 : ColourData = 12'hF8E;
20'b00000010100000010100 : ColourData = 12'hF8F;
20'b00000010110000010100 : ColourData = 12'hF8F;
20'b00000011000000010100 : ColourData = 12'hF8F;
20'b00000011010000010100 : ColourData = 12'hF9F;
20'b00000011100000010100 : ColourData = 12'hF9F;
20'b00000011110000010100 : ColourData = 12'h848;
20'b00000100000000010100 : ColourData = 12'h333;
20'b00000100010000010100 : ColourData = 12'h999;
20'b00000100100000010100 : ColourData = 12'h999;
20'b00000100110000010100 : ColourData = 12'h444;
20'b00000101000000010100 : ColourData = 12'h000;
20'b00000101010000010100 : ColourData = 12'h777;
20'b00000101100000010100 : ColourData = 12'h999;
20'b00000101110000010100 : ColourData = 12'h888;
20'b00000110000000010100 : ColourData = 12'h333;
20'b00000110010000010100 : ColourData = 12'h777;
20'b00000110100000010100 : ColourData = 12'h111;
20'b00000110110000010100 : ColourData = 12'h444;
20'b00000111000000010100 : ColourData = 12'h999;
20'b00000111010000010100 : ColourData = 12'h444;
20'b00000111100000010100 : ColourData = 12'h777;
20'b00000111110000010100 : ColourData = 12'hFFF;
20'b00000000000000010101 : ColourData = 12'h1F0;
20'b00000000010000010101 : ColourData = 12'h1F0;
20'b00000000100000010101 : ColourData = 12'h1F0;
20'b00000000110000010101 : ColourData = 12'h098;
20'b00000001000000010101 : ColourData = 12'h06B;
20'b00000001010000010101 : ColourData = 12'h013;
20'b00000001100000010101 : ColourData = 12'h000;
20'b00000001110000010101 : ColourData = 12'h975;
20'b00000010000000010101 : ColourData = 12'hF9E;
20'b00000010010000010101 : ColourData = 12'hF8F;
20'b00000010100000010101 : ColourData = 12'hF9F;
20'b00000010110000010101 : ColourData = 12'hF9F;
20'b00000011000000010101 : ColourData = 12'hF7E;
20'b00000011010000010101 : ColourData = 12'hF4B;
20'b00000011100000010101 : ColourData = 12'hF9F;
20'b00000011110000010101 : ColourData = 12'h848;
20'b00000100000000010101 : ColourData = 12'h233;
20'b00000100010000010101 : ColourData = 12'hB99;
20'b00000100100000010101 : ColourData = 12'hD99;
20'b00000100110000010101 : ColourData = 12'h877;
20'b00000101000000010101 : ColourData = 12'h666;
20'b00000101010000010101 : ColourData = 12'h888;
20'b00000101100000010101 : ColourData = 12'h999;
20'b00000101110000010101 : ColourData = 12'h999;
20'b00000110000000010101 : ColourData = 12'h777;
20'b00000110010000010101 : ColourData = 12'h888;
20'b00000110100000010101 : ColourData = 12'h666;
20'b00000110110000010101 : ColourData = 12'h977;
20'b00000111000000010101 : ColourData = 12'hE99;
20'b00000111010000010101 : ColourData = 12'h644;
20'b00000111100000010101 : ColourData = 12'h677;
20'b00000111110000010101 : ColourData = 12'hFFF;
20'b00000000000000010110 : ColourData = 12'h0C5;
20'b00000000010000010110 : ColourData = 12'h0C5;
20'b00000000100000010110 : ColourData = 12'h0C5;
20'b00000000110000010110 : ColourData = 12'h09D;
20'b00000001000000010110 : ColourData = 12'h09F;
20'b00000001010000010110 : ColourData = 12'h048;
20'b00000001100000010110 : ColourData = 12'h000;
20'b00000001110000010110 : ColourData = 12'h975;
20'b00000010000000010110 : ColourData = 12'hFAD;
20'b00000010010000010110 : ColourData = 12'hF8E;
20'b00000010100000010110 : ColourData = 12'hF7E;
20'b00000010110000010110 : ColourData = 12'hF8F;
20'b00000011000000010110 : ColourData = 12'hF7E;
20'b00000011010000010110 : ColourData = 12'hF4B;
20'b00000011100000010110 : ColourData = 12'hF9F;
20'b00000011110000010110 : ColourData = 12'h848;
20'b00000100000000010110 : ColourData = 12'h233;
20'b00000100010000010110 : ColourData = 12'hC99;
20'b00000100100000010110 : ColourData = 12'hF99;
20'b00000100110000010110 : ColourData = 12'hB99;
20'b00000101000000010110 : ColourData = 12'h788;
20'b00000101010000010110 : ColourData = 12'h888;
20'b00000101100000010110 : ColourData = 12'h888;
20'b00000101110000010110 : ColourData = 12'h777;
20'b00000110000000010110 : ColourData = 12'h999;
20'b00000110010000010110 : ColourData = 12'h888;
20'b00000110100000010110 : ColourData = 12'h777;
20'b00000110110000010110 : ColourData = 12'hC99;
20'b00000111000000010110 : ColourData = 12'hF99;
20'b00000111010000010110 : ColourData = 12'h744;
20'b00000111100000010110 : ColourData = 12'h677;
20'b00000111110000010110 : ColourData = 12'hFFF;
20'b00000000000000010111 : ColourData = 12'h08F;
20'b00000000010000010111 : ColourData = 12'h08F;
20'b00000000100000010111 : ColourData = 12'h08F;
20'b00000000110000010111 : ColourData = 12'h08F;
20'b00000001000000010111 : ColourData = 12'h08F;
20'b00000001010000010111 : ColourData = 12'h09F;
20'b00000001100000010111 : ColourData = 12'h025;
20'b00000001110000010111 : ColourData = 12'h974;
20'b00000010000000010111 : ColourData = 12'hFC9;
20'b00000010010000010111 : ColourData = 12'hF8D;
20'b00000010100000010111 : ColourData = 12'hF29;
20'b00000010110000010111 : ColourData = 12'hF8E;
20'b00000011000000010111 : ColourData = 12'hF9F;
20'b00000011010000010111 : ColourData = 12'hF8F;
20'b00000011100000010111 : ColourData = 12'hF9F;
20'b00000011110000010111 : ColourData = 12'h848;
20'b00000100000000010111 : ColourData = 12'h233;
20'b00000100010000010111 : ColourData = 12'hC99;
20'b00000100100000010111 : ColourData = 12'hF98;
20'b00000100110000010111 : ColourData = 12'hB99;
20'b00000101000000010111 : ColourData = 12'h333;
20'b00000101010000010111 : ColourData = 12'h777;
20'b00000101100000010111 : ColourData = 12'h888;
20'b00000101110000010111 : ColourData = 12'h111;
20'b00000110000000010111 : ColourData = 12'h888;
20'b00000110010000010111 : ColourData = 12'h777;
20'b00000110100000010111 : ColourData = 12'h000;
20'b00000110110000010111 : ColourData = 12'hB88;
20'b00000111000000010111 : ColourData = 12'hF99;
20'b00000111010000010111 : ColourData = 12'h744;
20'b00000111100000010111 : ColourData = 12'h667;
20'b00000111110000010111 : ColourData = 12'hFFF;
20'b00000000000000011000 : ColourData = 12'h09F;
20'b00000000010000011000 : ColourData = 12'h09F;
20'b00000000100000011000 : ColourData = 12'h09F;
20'b00000000110000011000 : ColourData = 12'h34F;
20'b00000001000000011000 : ColourData = 12'h42F;
20'b00000001010000011000 : ColourData = 12'h52F;
20'b00000001100000011000 : ColourData = 12'h105;
20'b00000001110000011000 : ColourData = 12'h974;
20'b00000010000000011000 : ColourData = 12'hFD9;
20'b00000010010000011000 : ColourData = 12'hFAA;
20'b00000010100000011000 : ColourData = 12'hF6D;
20'b00000010110000011000 : ColourData = 12'hF8F;
20'b00000011000000011000 : ColourData = 12'hF8F;
20'b00000011010000011000 : ColourData = 12'hF8F;
20'b00000011100000011000 : ColourData = 12'hF8F;
20'b00000011110000011000 : ColourData = 12'hD7D;
20'b00000100000000011000 : ColourData = 12'h646;
20'b00000100010000011000 : ColourData = 12'h655;
20'b00000100100000011000 : ColourData = 12'hB99;
20'b00000100110000011000 : ColourData = 12'hA99;
20'b00000101000000011000 : ColourData = 12'h222;
20'b00000101010000011000 : ColourData = 12'h222;
20'b00000101100000011000 : ColourData = 12'h222;
20'b00000101110000011000 : ColourData = 12'h000;
20'b00000110000000011000 : ColourData = 12'h222;
20'b00000110010000011000 : ColourData = 12'h111;
20'b00000110100000011000 : ColourData = 12'h000;
20'b00000110110000011000 : ColourData = 12'hA99;
20'b00000111000000011000 : ColourData = 12'h966;
20'b00000111010000011000 : ColourData = 12'h655;
20'b00000111100000011000 : ColourData = 12'hCCD;
20'b00000111110000011000 : ColourData = 12'hFFF;
20'b00000000000000011001 : ColourData = 12'h16F;
20'b00000000010000011001 : ColourData = 12'h16F;
20'b00000000100000011001 : ColourData = 12'h16F;
20'b00000000110000011001 : ColourData = 12'h42F;
20'b00000001000000011001 : ColourData = 12'h61F;
20'b00000001010000011001 : ColourData = 12'h40A;
20'b00000001100000011001 : ColourData = 12'h002;
20'b00000001110000011001 : ColourData = 12'h432;
20'b00000010000000011001 : ColourData = 12'hEB8;
20'b00000010010000011001 : ColourData = 12'hFC9;
20'b00000010100000011001 : ColourData = 12'hFBB;
20'b00000010110000011001 : ColourData = 12'hFAC;
20'b00000011000000011001 : ColourData = 12'hFAB;
20'b00000011010000011001 : ColourData = 12'hFAB;
20'b00000011100000011001 : ColourData = 12'hFAB;
20'b00000011110000011001 : ColourData = 12'hFBC;
20'b00000100000000011001 : ColourData = 12'hC89;
20'b00000100010000011001 : ColourData = 12'h554;
20'b00000100100000011001 : ColourData = 12'h777;
20'b00000100110000011001 : ColourData = 12'h999;
20'b00000101000000011001 : ColourData = 12'h666;
20'b00000101010000011001 : ColourData = 12'h444;
20'b00000101100000011001 : ColourData = 12'h444;
20'b00000101110000011001 : ColourData = 12'h444;
20'b00000110000000011001 : ColourData = 12'h444;
20'b00000110010000011001 : ColourData = 12'h444;
20'b00000110100000011001 : ColourData = 12'h555;
20'b00000110110000011001 : ColourData = 12'h666;
20'b00000111000000011001 : ColourData = 12'h555;
20'b00000111010000011001 : ColourData = 12'hBBB;
20'b00000111100000011001 : ColourData = 12'hFFF;
20'b00000111110000011001 : ColourData = 12'hFFF;
20'b00000000000000011010 : ColourData = 12'h61F;
20'b00000000010000011010 : ColourData = 12'h61F;
20'b00000000100000011010 : ColourData = 12'h61F;
20'b00000000110000011010 : ColourData = 12'h51F;
20'b00000001000000011010 : ColourData = 12'h51F;
20'b00000001010000011010 : ColourData = 12'h205;
20'b00000001100000011010 : ColourData = 12'h000;
20'b00000001110000011010 : ColourData = 12'h000;
20'b00000010000000011010 : ColourData = 12'hC97;
20'b00000010010000011010 : ColourData = 12'hEC8;
20'b00000010100000011010 : ColourData = 12'hEB8;
20'b00000010110000011010 : ColourData = 12'hEC8;
20'b00000011000000011010 : ColourData = 12'hEC8;
20'b00000011010000011010 : ColourData = 12'hEC8;
20'b00000011100000011010 : ColourData = 12'hEC8;
20'b00000011110000011010 : ColourData = 12'hEB8;
20'b00000100000000011010 : ColourData = 12'hFC8;
20'b00000100010000011010 : ColourData = 12'h864;
20'b00000100100000011010 : ColourData = 12'h555;
20'b00000100110000011010 : ColourData = 12'h999;
20'b00000101000000011010 : ColourData = 12'h999;
20'b00000101010000011010 : ColourData = 12'h999;
20'b00000101100000011010 : ColourData = 12'h999;
20'b00000101110000011010 : ColourData = 12'h999;
20'b00000110000000011010 : ColourData = 12'h999;
20'b00000110010000011010 : ColourData = 12'h999;
20'b00000110100000011010 : ColourData = 12'h999;
20'b00000110110000011010 : ColourData = 12'h444;
20'b00000111000000011010 : ColourData = 12'h555;
20'b00000111010000011010 : ColourData = 12'hFFF;
20'b00000111100000011010 : ColourData = 12'hFFF;
20'b00000111110000011010 : ColourData = 12'hFFF;
20'b00000000000000011011 : ColourData = 12'h51F;
20'b00000000010000011011 : ColourData = 12'h51F;
20'b00000000100000011011 : ColourData = 12'h51F;
20'b00000000110000011011 : ColourData = 12'hB9F;
20'b00000001000000011011 : ColourData = 12'h879;
20'b00000001010000011011 : ColourData = 12'h445;
20'b00000001100000011011 : ColourData = 12'h888;
20'b00000001110000011011 : ColourData = 12'h888;
20'b00000010000000011011 : ColourData = 12'h222;
20'b00000010010000011011 : ColourData = 12'h100;
20'b00000010100000011011 : ColourData = 12'h110;
20'b00000010110000011011 : ColourData = 12'h100;
20'b00000011000000011011 : ColourData = 12'h110;
20'b00000011010000011011 : ColourData = 12'h110;
20'b00000011100000011011 : ColourData = 12'h100;
20'b00000011110000011011 : ColourData = 12'h100;
20'b00000100000000011011 : ColourData = 12'h100;
20'b00000100010000011011 : ColourData = 12'h000;
20'b00000100100000011011 : ColourData = 12'h000;
20'b00000100110000011011 : ColourData = 12'h000;
20'b00000101000000011011 : ColourData = 12'h000;
20'b00000101010000011011 : ColourData = 12'h000;
20'b00000101100000011011 : ColourData = 12'h000;
20'b00000101110000011011 : ColourData = 12'h000;
20'b00000110000000011011 : ColourData = 12'h000;
20'b00000110010000011011 : ColourData = 12'h000;
20'b00000110100000011011 : ColourData = 12'h000;
20'b00000110110000011011 : ColourData = 12'h777;
20'b00000111000000011011 : ColourData = 12'hEEE;
20'b00000111010000011011 : ColourData = 12'hFFF;
20'b00000111100000011011 : ColourData = 12'hFFF;
20'b00000111110000011011 : ColourData = 12'hFFF;
20'b00000000000000011100 : ColourData = 12'h73E;
20'b00000000010000011100 : ColourData = 12'h74F;
20'b00000000100000011100 : ColourData = 12'h74E;
20'b00000000110000011100 : ColourData = 12'hEDF;
20'b00000001000000011100 : ColourData = 12'h9A9;
20'b00000001010000011100 : ColourData = 12'h555;
20'b00000001100000011100 : ColourData = 12'h999;
20'b00000001110000011100 : ColourData = 12'h666;
20'b00000010000000011100 : ColourData = 12'h011;
20'b00000010010000011100 : ColourData = 12'h666;
20'b00000010100000011100 : ColourData = 12'h111;
20'b00000010110000011100 : ColourData = 12'h444;
20'b00000011000000011100 : ColourData = 12'h333;
20'b00000011010000011100 : ColourData = 12'h011;
20'b00000011100000011100 : ColourData = 12'h888;
20'b00000011110000011100 : ColourData = 12'h888;
20'b00000100000000011100 : ColourData = 12'h888;
20'b00000100010000011100 : ColourData = 12'h888;
20'b00000100100000011100 : ColourData = 12'h222;
20'b00000100110000011100 : ColourData = 12'h222;
20'b00000101000000011100 : ColourData = 12'h555;
20'b00000101010000011100 : ColourData = 12'h000;
20'b00000101100000011100 : ColourData = 12'h666;
20'b00000101110000011100 : ColourData = 12'h000;
20'b00000110000000011100 : ColourData = 12'h444;
20'b00000110010000011100 : ColourData = 12'h333;
20'b00000110100000011100 : ColourData = 12'h000;
20'b00000110110000011100 : ColourData = 12'hCCC;
20'b00000111000000011100 : ColourData = 12'hFFF;
20'b00000111010000011100 : ColourData = 12'hFFF;
20'b00000111100000011100 : ColourData = 12'hFFF;
20'b00000111110000011100 : ColourData = 12'hFFF;
20'b00000000000000011101 : ColourData = 12'hFFF;
20'b00000000010000011101 : ColourData = 12'hFFF;
20'b00000000100000011101 : ColourData = 12'hFFF;
20'b00000000110000011101 : ColourData = 12'hFFF;
20'b00000001000000011101 : ColourData = 12'h999;
20'b00000001010000011101 : ColourData = 12'h444;
20'b00000001100000011101 : ColourData = 12'h888;
20'b00000001110000011101 : ColourData = 12'h555;
20'b00000010000000011101 : ColourData = 12'h777;
20'b00000010010000011101 : ColourData = 12'hCCD;
20'b00000010100000011101 : ColourData = 12'h222;
20'b00000010110000011101 : ColourData = 12'h777;
20'b00000011000000011101 : ColourData = 12'h666;
20'b00000011010000011101 : ColourData = 12'h444;
20'b00000011100000011101 : ColourData = 12'hFFF;
20'b00000011110000011101 : ColourData = 12'hFFF;
20'b00000100000000011101 : ColourData = 12'hFFF;
20'b00000100010000011101 : ColourData = 12'hFFF;
20'b00000100100000011101 : ColourData = 12'h666;
20'b00000100110000011101 : ColourData = 12'h556;
20'b00000101000000011101 : ColourData = 12'h888;
20'b00000101010000011101 : ColourData = 12'h111;
20'b00000101100000011101 : ColourData = 12'hCCC;
20'b00000101110000011101 : ColourData = 12'h334;
20'b00000110000000011101 : ColourData = 12'h888;
20'b00000110010000011101 : ColourData = 12'h666;
20'b00000110100000011101 : ColourData = 12'h334;
20'b00000110110000011101 : ColourData = 12'hFFF;
20'b00000111000000011101 : ColourData = 12'hFFF;
20'b00000111010000011101 : ColourData = 12'hFFF;
20'b00000111100000011101 : ColourData = 12'hFFF;
20'b00000111110000011101 : ColourData = 12'hFFF;
20'b00000000000000011110 : ColourData = 12'hFFF;
20'b00000000010000011110 : ColourData = 12'hFFF;
20'b00000000100000011110 : ColourData = 12'hFFF;
20'b00000000110000011110 : ColourData = 12'hFFF;
20'b00000001000000011110 : ColourData = 12'h999;
20'b00000001010000011110 : ColourData = 12'h000;
20'b00000001100000011110 : ColourData = 12'h000;
20'b00000001110000011110 : ColourData = 12'h000;
20'b00000010000000011110 : ColourData = 12'hCCC;
20'b00000010010000011110 : ColourData = 12'hFFF;
20'b00000010100000011110 : ColourData = 12'h111;
20'b00000010110000011110 : ColourData = 12'h000;
20'b00000011000000011110 : ColourData = 12'h333;
20'b00000011010000011110 : ColourData = 12'hEEE;
20'b00000011100000011110 : ColourData = 12'hFFF;
20'b00000011110000011110 : ColourData = 12'hFFF;
20'b00000100000000011110 : ColourData = 12'hFFF;
20'b00000100010000011110 : ColourData = 12'hFFF;
20'b00000100100000011110 : ColourData = 12'hEEE;
20'b00000100110000011110 : ColourData = 12'h555;
20'b00000101000000011110 : ColourData = 12'h000;
20'b00000101010000011110 : ColourData = 12'h000;
20'b00000101100000011110 : ColourData = 12'hDDD;
20'b00000101110000011110 : ColourData = 12'hEEE;
20'b00000110000000011110 : ColourData = 12'h111;
20'b00000110010000011110 : ColourData = 12'h333;
20'b00000110100000011110 : ColourData = 12'hEEE;
20'b00000110110000011110 : ColourData = 12'hFFF;
20'b00000111000000011110 : ColourData = 12'hFFF;
20'b00000111010000011110 : ColourData = 12'hFFF;
20'b00000111100000011110 : ColourData = 12'hFFF;
20'b00000111110000011110 : ColourData = 12'hFFF;
20'b00000000000000011111 : ColourData = 12'hFFF;
20'b00000000010000011111 : ColourData = 12'hFFF;
20'b00000000100000011111 : ColourData = 12'hFFF;
20'b00000000110000011111 : ColourData = 12'hFFF;
20'b00000001000000011111 : ColourData = 12'hEEE;
20'b00000001010000011111 : ColourData = 12'hBBB;
20'b00000001100000011111 : ColourData = 12'hBBB;
20'b00000001110000011111 : ColourData = 12'hCCC;
20'b00000010000000011111 : ColourData = 12'hEFF;
20'b00000010010000011111 : ColourData = 12'hFFF;
20'b00000010100000011111 : ColourData = 12'hCCC;
20'b00000010110000011111 : ColourData = 12'hBBB;
20'b00000011000000011111 : ColourData = 12'hCCD;
20'b00000011010000011111 : ColourData = 12'hFFF;
20'b00000011100000011111 : ColourData = 12'hFFF;
20'b00000011110000011111 : ColourData = 12'hFFF;
20'b00000100000000011111 : ColourData = 12'hFFF;
20'b00000100010000011111 : ColourData = 12'hFFF;
20'b00000100100000011111 : ColourData = 12'hFFF;
20'b00000100110000011111 : ColourData = 12'hDDD;
20'b00000101000000011111 : ColourData = 12'hBCC;
20'b00000101010000011111 : ColourData = 12'hCCC;
20'b00000101100000011111 : ColourData = 12'hFFF;
20'b00000101110000011111 : ColourData = 12'hFFF;
20'b00000110000000011111 : ColourData = 12'hCCC;
20'b00000110010000011111 : ColourData = 12'hDDD;
20'b00000110100000011111 : ColourData = 12'hFFF;
20'b00000110110000011111 : ColourData = 12'hFFF;
20'b00000111000000011111 : ColourData = 12'hFFF;
20'b00000111010000011111 : ColourData = 12'hFFF;
20'b00000111100000011111 : ColourData = 12'hFFF;
20'b00000111110000011111 : ColourData = 12'hFFF;



default: ColourData = 12'h000;

endcase
end

endmodule
