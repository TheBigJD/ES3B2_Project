module VGA_Draw(
    input Master_Clock_In, Reset_N_In,
    input Disp_Ena_In,
    input [9:0] Val_Col_In, Val_Row_In,
    
    input Up, Down, Left, Right, Fire,
    
    input LevelSwitch_1, LevelSwitch_0,
    input ColourSwitch_1,
    input MoveSpeed_1, MoveSpeed_0,
    
	output reg [7:0] CoinValue = 8'd0,
	output reg debug_led = 1'b0, // test LED for debugging
	
	output reg [3:0] Red   = 4'h0, 
	output reg [3:0] Blue  = 4'h0, 
    output reg [3:0] Green = 4'h0
);

parameter Pixels_Horiz = 640; //Num of Pixels in X axis
parameter Pixels_Vert  = 480; //Num of Pixels in Y axis

parameter EdgeWidth = 0;

parameter [2:0] Up_Direction      = 3'b100;	
parameter [2:0] Down_Direction    = 3'b001;	
parameter [2:0] Left_Direction    = 3'b010;	
parameter [2:0] Right_Direction   = 3'b011;	

parameter TankWidth   = 24;

reg [2:0] MoveSpeed = 3'b1;
	
parameter [3:0] BulletWidth = 4'd10; // Square bullet
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

reg [9:0] PrevX, PrevY = 10'b0;

reg [2:0] PrevDirection = 3'b00;	

reg [9:0] Tank1_xPos = 10'd4;
reg [9:0] Tank1_yPos = 10'd4;	
	
reg [9:0] xDivPos, yDivPos= 10'b0;	
	
reg [9:0] Tank_xDivPos_1, Tank_yDivPos_1;
reg [9:0] Tank_xDivPos_2, Tank_yDivPos_2;
reg [9:0] Tank1_xPos2_Holder, Tank1_yPos2_Holder;

reg [0:79] TankArray_1 = 80'b0;
reg [3:0] TankArray_X_1 = 4'b0;
reg TankArray_1_0, TankArray_1_1, TankArray_1_2, TankArray_1_3;

reg [0:79] TankArray_2 = 80'b0;
reg [3:0] TankArray_X_2 = 4'b0;
reg TankArray_2_0, TankArray_2_1, TankArray_2_2, TankArray_2_3;

reg [0:79] TankArray_3 = 80'b0;
reg [3:0] TankArray_X_3 = 4'b0;
reg TankArray_3_0, TankArray_3_1, TankArray_3_2, TankArray_3_3;

reg [0:79] TankArray_4 = 80'b0;
reg [3:0] TankArray_X_4 = 4'b0;
reg TankArray_4_0, TankArray_4_1, TankArray_4_2, TankArray_4_3;



///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Instantiating colour inputs

wire [11:0] Colour_Data_Background;
//Bottle M4 (.Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Background));

reg [9:0] Tank_XInput, Tank_YInput = 10'b0;	
wire [11:0] Colour_Data_Tank;
TankImage M5 (.Master_Clock_In(Master_Clock_In), .xInput(Tank_XInput), .yInput(Tank_YInput), .ColourData(Colour_Data_Tank));

wire [11:0] Colour_Data_Brick;
Brick_Block M6( .Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Brick));

wire [11:0] Colour_Data_Nyan;
MysteryImage M7( .Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Nyan));

wire [11:0] Colour_Data_Solid_Block;
Solid_block M8( .Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Solid_Block));
	
wire [11:0] Colour_Data_Coin;
Coin_Image M9( .Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In), .yInput(Val_Col_In), .ColourData(Colour_Data_Coin));

reg [9:0] Bullet_XInput_1, Bullet_YInput_1 = 10'd16; // TODO does this only set Yinput to d16?
wire [11:0] Colour_Data_Bullet;
Bullet M10( .Master_Clock_In(Master_Clock_In), .xInput(Val_Row_In - Bullet_XInput_1 - BulletWidth/2), .yInput(Val_Col_In - Bullet_YInput_1 - BulletWidth/2), .ColourData(Colour_Data_Bullet));


	
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Bullets?


reg Bullet_Fired_prev_1 = 1'b0;
reg Bullet_Fired_prev_2 = 1'b0;
reg Bullet_Fired_1		= 1'b0;
reg [2:0] Bullet_Dir_1  = 2'b000;

reg [5:0] Bullet_ClockDiv = 6'b0;
reg [5:0] Bullet_ClockCounter = 6'd30;
	// Note - these are coded differently to the tank bounding boxes. Tanks are done at each corner, whereas this is done
	//		at the centre only
	
//reg [0:79] BulletArray_1 = 80'b0;
reg [3:0] BulletArray_X = 4'b0;
reg [0:79] BulletArrayData_Y = 80'b0;
reg BulletArrayData_X_0, BulletArrayData_X_1, BulletArrayData_X_2, BulletArrayData_X_3;

reg [9:0] Bullet_xDivPos_1, Bullet_yDivPos_1 = 10'b0;
	
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
	
reg [0:79] MapArray [0:14];
reg [0:79] MapArrayData_Y = 80'b0;
reg [3:0]  MapArray_X = 4'b0;
reg MapArrayData_X_3, MapArrayData_X_2, MapArrayData_X_1, MapArrayData_X_0;



always @(posedge Master_Clock_In)	
	begin
		if (Reset_N_In == 0)
			begin
                Red   = 4'h0;     
                Blue  = 4'h0;
                Green = 4'h0;
                    
                Bullet_Fired_1 = 1'b0; // TODO defined twice - should this be reset on every posedge? 
                Bullet_XInput_1 = 10'd16; 
                Bullet_YInput_1 = 10'd16;
                Tank1_xPos = 10'd5;
                Tank1_yPos = 10'd5;
                CoinValue = 8'd0;
				
				case ({LevelSwitch_1, LevelSwitch_0})
					3: begin
						MapArray[ 0] = 80'b0001_0001_0001_0001_0001_0001_0001_0001_0000_0001_0001_0001_0001_0001_0000_0001_0001_0001_0001_0001;
                        MapArray[ 1] = 80'b0001_0010_0000_0000_0000_0010_0010_0010_0000_0010_0010_0010_0010_0010_0000_0000_0010_0000_0101_0001;
                        MapArray[ 2] = 80'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000;
                        MapArray[ 3] = 80'b0001_0000_0000_0010_0010_0010_0000_0000_0001_0010_0001_0000_0000_0010_0000_0001_0001_0001_0000_0001;
                        MapArray[ 4] = 80'b0001_0000_0010_0010_0101_0000_0000_0001_0001_0101_0001_0001_0000_0000_0000_0000_0000_0000_0000_0001;
                        MapArray[ 5] = 80'b0001_0000_0010_0001_0101_0000_0000_0010_0101_0101_0101_0010_0000_0010_0001_0010_0010_0010_0001_0001;
                        MapArray[ 6] = 80'b0001_0000_0000_0001_0001_0001_0000_0010_0101_0101_0101_0000_0000_0001_0001_0101_0101_0101_0001_0001;
                        MapArray[ 7] = 80'b0001_0000_0000_0000_0000_0000_0000_0001_0001_0101_0001_0001_0000_0010_0001_0010_0010_0010_0001_0001;
                        MapArray[ 8] = 80'b0000_0000_0001_0000_0010_0000_0000_0000_0001_0010_0001_0010_0000_0000_0000_0000_0000_0000_0000_0000;
                        MapArray[ 9] = 80'b0001_0000_0001_0000_0001_0000_0001_0000_0010_0000_0000_0010_0000_0010_0010_0001_0001_0001_0010_0001;
                        MapArray[10] = 80'b0001_0000_0001_0101_0001_0000_0000_0000_0010_0000_0000_0010_0000_0001_0010_0101_0101_0101_0010_0001;
                        MapArray[11] = 80'b0001_0000_0000_0001_0000_0000_0000_0000_0010_0101_0010_0001_0000_0010_0010_0001_0001_0001_0010_0001;
                        MapArray[12] = 80'b0001_0010_0000_0000_0000_0001_0001_0000_0001_0010_0010_0000_0000_0000_0000_0000_0000_0000_0000_0001;
                        MapArray[13] = 80'b0001_0010_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0010_0000_0000_0101_0001;
                        MapArray[14] = 80'b0001_0001_0001_0001_0001_0001_0001_0001_0000_0001_0001_0001_0001_0001_0000_0001_0001_0001_0001_0001;
	

					end
						
					2: begin // Pacman level
						MapArray[ 0] = 80'h11111111111111111111;
						MapArray[ 1] = 80'h13331333333333313331;
						MapArray[ 2] = 80'h13131331133113313131;
						MapArray[ 3] = 80'h13133333333333333131;
						MapArray[ 4] = 80'h13113113133131131131;
						MapArray[ 5] = 80'h13313333133133331331;
						MapArray[ 6] = 80'h03311313333331311330;
						MapArray[ 7] = 80'h03333311111111333330;
						MapArray[ 8] = 80'h13313333333333331331;
						MapArray[ 9] = 80'h11311131111113111311;
						MapArray[10] = 80'h13333133333333133331;
						MapArray[11] = 80'h13113331111113331131;
						MapArray[12] = 80'h13113131111113131131;
						MapArray[13] = 80'h13333133333333133331;
						MapArray[14] = 80'h11111111111111111111;
					end
					
				    1: begin
				        MapArray[ 0] = 80'b0001_0001_0001_0000_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0000_0001_0001_0001;
                        MapArray[ 1] = 80'b0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001;
                        MapArray[ 2] = 80'b0001_0011_0001_0001_0001_0011_0010_0010_0011_0000_0000_0011_0010_0010_0011_0001_0001_0001_0011_0001;
                        MapArray[ 3] = 80'b0001_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0001;
                        MapArray[ 4] = 80'b0001_0000_0010_0010_0010_0000_0010_0000_0001_0001_0001_0001_0000_0010_0000_0010_0010_0010_0000_0001;
                        MapArray[ 5] = 80'b0001_0000_0000_0000_0000_0000_0010_0000_0000_0010_0010_0000_0000_0010_0000_0000_0000_0000_0000_0001;
                        MapArray[ 6] = 80'b0001_0000_0001_0000_0000_0010_0010_0000_0000_0010_0010_0000_0000_0010_0010_0000_0000_0001_0000_0001;
                        MapArray[ 7] = 80'b0000_0000_0001_0011_0010_0011_0011_0010_0011_0010_0010_0011_0010_0011_0011_0010_0011_0001_0000_0000;
                        MapArray[ 8] = 80'b0001_0000_0001_0000_0000_0010_0010_0000_0000_0010_0010_0000_0000_0010_0010_0000_0000_0001_0000_0001;
                        MapArray[ 9] = 80'b0001_0000_0000_0000_0000_0000_0010_0000_0000_0010_0010_0000_0000_0010_0000_0000_0000_0000_0000_0001;
                        MapArray[10] = 80'b0001_0000_0010_0010_0010_0000_0010_0000_0001_0001_0001_0001_0000_0010_0000_0010_0010_0010_0000_0001;
                        MapArray[11] = 80'b0001_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0001;
                        MapArray[12] = 80'b0001_0011_0001_0001_0001_0011_0010_0010_0011_0000_0000_0011_0010_0010_0011_0001_0001_0001_0011_0001;
                        MapArray[13] = 80'b0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001;
                        MapArray[14] = 80'b0001_0001_0001_0000_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0001_0000_0001_0001_0001;
                    end
				    
				    
				    0: begin//coin
                        MapArray[ 0] = 80'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
                        MapArray[ 1] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                        MapArray[ 2] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                        MapArray[ 3] = 80'b0000_0010_0010_0010_0010_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0010_0010_0010_0010_0000;
                        MapArray[ 4] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                        MapArray[ 5] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0010_0010_0010_0011_0010_0010_0011_0010_0011_0011_0000;
                        MapArray[ 6] = 80'b0000_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0000;
                        MapArray[ 7] = 80'b0000_0010_0010_0010_0010_0010_0011_0010_0010_0010_0010_0010_0010_0011_0010_0010_0010_0010_0010_0000;
                        MapArray[ 8] = 80'b0000_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0011_0000;
                        MapArray[ 9] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0010_0010_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                        MapArray[10] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                        MapArray[11] = 80'b0000_0010_0010_0010_0010_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0010_0010_0010_0010_0000;
                        MapArray[12] = 80'b0000_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0010_0011_0011_0011_0011_0010_0011_0011_0000;
                        MapArray[13] = 80'b0000_0010_0011_0010_0011_0010_0010_0011_0010_0011_0011_0010_0011_0010_0010_0011_0010_0011_0010_0000;
                        MapArray[14] = 80'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        			end
                    
                endcase
			end
		else 
			begin
			// Need control for map choice here
            if (Disp_Ena_In == 0)
                begin
                    Red 	= {4{1'b0}};
                    Blue 	= {4{1'b0}};
                    Green 	= {4{1'b0}};
                end
        
            else
                begin
                    if ((Val_Col_In <= Pixels_Vert) & (Val_Row_In <= Pixels_Horiz)) 
                        begin

////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                            //do not delete this. or i kill you.
                            // this is the bit that takes the x/y coordinates and shuffles them into the 20by15 array
                            // This will give the data for essentially 'What should we do with the tank at this point?
                            // We need to observe points at (x, y), (x+w, y), (x,y+w), (x+w, y+w) and make sure that these points
                            //      that the tank movement is limited if it reaches a point where the tank cant move through.
                            // This will allow the basis for the bullets too. If it hits a breakable block, we can change the reg's
                            //      value at this point to 4'h0, and the tank will behave differently than it would if it was 4'h2.
                            if ((Val_Col_In == Pixels_Vert) & (Val_Row_In == Pixels_Horiz))
                                begin
							// There might be a better way of ordering these values - overwriting might make an impact
							//	on gameplay
////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////
									//Bullet controls

									//Rising edge of 'Fire' button input
									
                                    Bullet_Fired_prev_2 = Bullet_Fired_prev_1;
                                    Bullet_Fired_prev_1 = Fire; 
                                    
                                    if ((Fire == 1'b1) & (Bullet_Fired_prev_2 == 1'b0) & (Bullet_Fired_1 == 0)) // Create new bullet as no other bullets currently on screen
                                    //if ((Bullet_Fired_prev_1 == 0) & (Fire == 1))
                                        begin
                                            Bullet_Fired_1   = 1'b1; // Bullet is now enabled
                                            Bullet_Dir_1    = PrevDirection; // Use same direction as movement of tank for bullet
                                            
                                            case (Bullet_Dir_1) // Define initial bullet position depending on direction
                                                Up_Direction:
                                                    begin
                                                        Bullet_XInput_1 = Tank1_xPos + (BulletWidth + 3);
                                                        Bullet_YInput_1 = Tank1_yPos - (BulletWidth + 3);
                                                    end
                                                    
                                                Down_Direction:
                                                    begin
                                                        Bullet_XInput_1 = Tank1_xPos + (BulletWidth + 3);
                                                        Bullet_YInput_1 = Tank1_yPos + (BulletWidth + 3) + TankWidth;
                                                    end
                                                    
                                                Left_Direction:
                                                    begin
                                                        Bullet_XInput_1 = Tank1_xPos - (BulletWidth + 3);
                                                        Bullet_YInput_1 = Tank1_yPos + (BulletWidth + 3);
                                                    end
                                                    
                                                Right_Direction:
                                                    begin
                                                        Bullet_XInput_1 = Tank1_xPos + (BulletWidth + 3) + TankWidth;
                                                        Bullet_YInput_1 = Tank1_yPos - (BulletWidth + 3) + TankWidth;
                                                    end
                                                    
                                                default: Bullet_Fired_1 = 1'b0; //TODO is this the correct place to set Bullet_fired_1 off? presumably Bullet_Dir_1 only gets 4 possible direction inputs; all are covered above
                                            endcase
                                        end
                                        
                                    else if (Bullet_Fired_1 == 1) // continue moving bullet across screen
                                        begin
                                            Bullet_xDivPos_1 = (Bullet_XInput_1[9:5])%20;
                                            Bullet_yDivPos_1 = (Bullet_YInput_1[9:5])%15;
                                            
                                            BulletArrayData_Y   = MapArray[Bullet_yDivPos_1]; // 
                                            BulletArrayData_X_3 = BulletArrayData_Y[4* (Bullet_xDivPos_1)];
                                            BulletArrayData_X_2 = BulletArrayData_Y[4* (Bullet_xDivPos_1) + 1];
                                            BulletArrayData_X_1 = BulletArrayData_Y[4* (Bullet_xDivPos_1) + 2];
                                            BulletArrayData_X_0 = BulletArrayData_Y[4* (Bullet_xDivPos_1) + 3];
                                            
                                            BulletArray_X = {BulletArrayData_X_3, BulletArrayData_X_2, BulletArrayData_X_1, BulletArrayData_X_0 };
                                            
                                            //Define what happens when bullet hits edges of screen
                                            if ((Bullet_XInput_1 <= BulletWidth) | (Bullet_YInput_1 <= BulletWidth) | (Bullet_XInput_1 >= Pixels_Horiz - BulletWidth) | (Bullet_YInput_1 >= Pixels_Vert - BulletWidth))
                                                begin
                                                    Bullet_XInput_1 = 10'd16; // Reset bullet position to default X and Y
                                                    Bullet_YInput_1 = 10'd16;
                                                    Bullet_Fired_1 	=  1'b0; // Stop firing bullet
                                                end
                                            
                                            // if hit tank                                            
                                            if ((BulletArray_X == 1) | (BulletArray_X == 2)) // TODO When is BulletArray_X either of these values?
                                                begin
                                                    Bullet_XInput_1 = 10'd16; // Reset bullet position to default X and Y
                                                    Bullet_YInput_1 = 10'd16;
                                                    Bullet_Fired_1 	=  1'b0; // Stop firing bullet
                                    
                                                    if (BulletArray_X == 2)
                                                        begin
                                                            MapArray[Bullet_yDivPos_1][4 * Bullet_xDivPos_1	   ] = 1'b0;	
                                                            MapArray[Bullet_yDivPos_1][4 * Bullet_xDivPos_1 + 1] = 1'b0;
                                                            MapArray[Bullet_yDivPos_1][4 * Bullet_xDivPos_1 + 2] = 1'b0;
                                                            MapArray[Bullet_yDivPos_1][4 * Bullet_xDivPos_1 + 3] = 1'b0;
                                                        end
                                                end
                                                
                                            else if ((BulletArray_X == 0) | (BulletArray_X == 3))  
                                           
                                                begin
                                                    case (Bullet_Dir_1)
                                                    
                                                        Up_Direction    : Bullet_YInput_1 = Bullet_YInput_1 - 5;
                                                        Down_Direction  : Bullet_YInput_1 = Bullet_YInput_1 + 5;
                                                        Left_Direction  : Bullet_XInput_1 = Bullet_XInput_1 - 5;
                                                        Right_Direction : Bullet_XInput_1 = Bullet_XInput_1 + 5;
                                                        default: Bullet_Fired_1 = 1'b0;
                                                    endcase	
                                                end
                                            else
                                                begin
                                                    Bullet_XInput_1 = 10'd16; // Reset bullet position to default X and Y
                                                    Bullet_YInput_1 = 10'd16;
                                                    Bullet_Fired_1 	=  1'b0; // Stop firing bullet
                                                end
                                        end
                                    else
                                        begin
                                            Bullet_XInput_1 = 10'b0;
                                            Bullet_YInput_1 = 10'b0;
                                            Bullet_Fired_1 	= 1'b0;
                                        end
////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                                    // If y-coordinate is at screen limit, move to other side of screen
//                                    if (Tank1_yPos <= EdgeWidth)
//                                        begin
//                                            Tank1_yPos = Pixels_Vert - TankWidth - 1;
//                                        end
//                                    else if (Tank1_yPos >= Pixels_Vert - TankWidth - EdgeWidth)
//                                        begin
//                                            Tank1_yPos = 10'd3;
//                                        end
//                                    //if x-coordinate is at screen limit, move to other side of screen
//                                    else if (Tank1_xPos <= EdgeWidth) // TODO add else?
//                                        begin
//                                            Tank1_xPos = Pixels_Horiz - TankWidth - 1;
//                                        end
//                                    else if (Tank1_xPos >= Pixels_Horiz - TankWidth - EdgeWidth)
//                                        begin
//                                            Tank1_xPos = 10'd3;
//                                        end
////////////////////////////////////////////////////////////////////////////////////////////////////////////////                    
////////////////////////////////////////////////////////////////////////////////////////////////////////////////                    
                                    //Setting Bounding boxes for tank control. Looking for box state at x and y positions
                                    Tank_xDivPos_1 = Tank1_xPos[9:5]%20;
                                    Tank_yDivPos_1 = Tank1_yPos[9:5]%15;
                                    
									Tank1_xPos2_Holder = Tank1_xPos + TankWidth;
									Tank1_yPos2_Holder = Tank1_xPos2_Holder[9:5]%20;
                                    Tank_yDivPos_2 = Tank1_yPos2_Holder[9:5]%15;
                                   
//////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////  
                                    //Top left
                                    TankArray_1   = MapArray[Tank_yDivPos_1];// This is the array for the map containing the 'bottom left#' of the tank
                                    TankArray_1_3 = TankArray_1[4*Tank_xDivPos_1  ];// This is bit 3 of [3:0] of the current position's status.
                                    TankArray_1_2 = TankArray_1[4*Tank_xDivPos_1+1];// This is bit 2 of [3:0] of the current position's status.
                                    TankArray_1_1 = TankArray_1[4*Tank_xDivPos_1+2];// This is bit 1 of [3:0] of the current position's status.v
                                    TankArray_1_0 = TankArray_1[4*Tank_xDivPos_1+3];// This is bit 0 of [3:0] of the current position's status.
									
                                    TankArray_X_1 = {TankArray_1_3, TankArray_1_2, TankArray_1_1, TankArray_1_0};
									//This then returns the state of the box for the bottom-left point of the tank, allowing for the game logic to perform functions depending
									//		on the position of the tank.
									
									// The same logic repeats for each corner of the tank.

                                    //Top right
                                    TankArray_2   = MapArray[Tank_yDivPos_1];
                                    TankArray_2_3 = TankArray_2[4*(Tank_xDivPos_2 )  ];
                                    TankArray_2_2 = TankArray_2[4*(Tank_xDivPos_2 )+1];
                                    TankArray_2_1 = TankArray_2[4*(Tank_xDivPos_2 )+2];
                                    TankArray_2_0 = TankArray_2[4*(Tank_xDivPos_2 )+3];
                                    TankArray_X_2 = {TankArray_2_3, TankArray_2_2, TankArray_2_1, TankArray_2_0}; 
									
                                    //Bottom left
                                    TankArray_3   = MapArray[Tank_yDivPos_2 ];
                                    TankArray_3_3 = TankArray_3[4*(Tank_xDivPos_1)  ];
                                    TankArray_3_2 = TankArray_3[4*(Tank_xDivPos_1)+1];
                                    TankArray_3_1 = TankArray_3[4*(Tank_xDivPos_1)+2];
                                    TankArray_3_0 = TankArray_3[4*(Tank_xDivPos_1)+3];
                                    TankArray_X_3 = {TankArray_3_3, TankArray_3_2, TankArray_3_1, TankArray_3_0};   
									
                                    //Bottom right
                                    TankArray_4   = MapArray[Tank_yDivPos_2 ];
                                    TankArray_4_3 = TankArray_4[4*(Tank_xDivPos_2 )  ];
                                    TankArray_4_2 = TankArray_4[4*(Tank_xDivPos_2 )+1];
                                    TankArray_4_1 = TankArray_4[4*(Tank_xDivPos_2 )+2];
                                    TankArray_4_0 = TankArray_4[4*(Tank_xDivPos_2 )+3];
                                    TankArray_X_4 = {TankArray_4_3, TankArray_4_2, TankArray_4_1, TankArray_4_0};   
									
///////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////  
                                    // If y-coordinate is at screen limit, move to other side of screen
                                    if (Tank1_yPos <= EdgeWidth)
                                        begin
                                            Tank1_yPos = Pixels_Vert - TankWidth - 3;
                                        end
                                    else if (Tank1_yPos >= Pixels_Vert - TankWidth - EdgeWidth)
                                        begin
                                            Tank1_yPos = 3;
                                        end

                                    //if x-coordinate is at screen limit, move to other side of screen
                                    else if (Tank1_xPos <= EdgeWidth)
                                        begin
                                            Tank1_xPos = Pixels_Horiz - TankWidth - 3;
                                        end
                                    else if (Tank1_xPos >= Pixels_Horiz - TankWidth - EdgeWidth)
                                        begin
                                            Tank1_xPos = 3;
                                        end
///////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////       
     
                                    //If bottom edges are in boundary
									else if (((TankArray_X_3 == 1) | (TankArray_X_3 == 2)) & ((TankArray_X_4 == 1) | (TankArray_X_4 == 2)))
                                        begin
                                            Tank1_yPos = Tank1_yPos - 1;
                                        end
												
                                    //If left edges are in boundary
								    else if (((TankArray_X_1 == 1) | (TankArray_X_1 == 2)) & ((TankArray_X_3 == 1) | (TankArray_X_3 == 2)))
                                        begin
                                            Tank1_xPos = Tank1_xPos + 1;
                                        end
												
                                    //if top edges are in boundary
                                    else if (((TankArray_X_1 == 1) | (TankArray_X_1 == 2)) & ((TankArray_X_2 == 1) | (TankArray_X_2 == 2)))
                                        begin
                                            Tank1_yPos = Tank1_yPos + 1;
                                        end
                                                    
                                    // if right edges are in boundary
                                    else if (((TankArray_X_2 == 1) | (TankArray_X_2 == 2)) & ((TankArray_X_4 == 1) | (TankArray_X_4 == 2)))
                                        begin
                                            Tank1_xPos = Tank1_xPos - 1;            
                                        end 
///////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////                                          
									// if top left is in boundary
									else if ((TankArray_X_1 == 1) | (TankArray_X_1 == 2))
										begin
											Tank1_yPos = Tank1_yPos + 1;
											Tank1_xPos = Tank1_xPos + 1;
										end
									// if top right is in boundary	
									else if ((TankArray_X_2 == 1) | (TankArray_X_2 == 2))
										begin
											Tank1_yPos = Tank1_yPos + 1;
											Tank1_xPos = Tank1_xPos - 1;
										end	
									// if bottom left is in boundary	
									else if ((TankArray_X_3 == 1) | (TankArray_X_3 == 2))
										begin
											Tank1_yPos = Tank1_yPos - 1;
											Tank1_xPos = Tank1_xPos + 1;
										end
									// if bottom right is in boundary	
									else if ((TankArray_X_4 == 1) | (TankArray_X_4 == 2))
										begin
											Tank1_yPos = Tank1_yPos - 1;
											Tank1_xPos = Tank1_xPos - 1;
										end	

///////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
									else if (TankArray_X_1 == 3)
										begin
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_1   ] = 1'b0;	
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_1+ 1] = 1'b0;	
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_1+ 2] = 1'b0;
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_1+ 3] = 1'b0;
											
											CoinValue = CoinValue + 1;	
											
										end
								
 									else if (TankArray_X_2 == 3)
										begin
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_2	 ]   = 1'b0;	
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_2 + 1] = 1'b0;
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_2 + 2] = 1'b0;
											MapArray[Tank_yDivPos_1][4 * Tank_xDivPos_2 + 3] = 1'b0;
											
											CoinValue = CoinValue + 1;
											
										end
								
 									else if (TankArray_X_3 == 3)
										begin
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_1   ] = 1'b0;	
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_1+ 1] = 1'b0;
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_1+ 2] = 1'b0;
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_1+ 3] = 1'b0;
											
											CoinValue = CoinValue + 1;
											
										end
								
 									else if (TankArray_X_4 == 3)
										begin
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_2   ] = 1'b0;	
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_2+ 1] = 1'b0;
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_2+ 2] = 1'b0;
											MapArray[Tank_yDivPos_2][4 * Tank_xDivPos_2+ 3] = 1'b0;
											
											CoinValue = CoinValue + 1;
											
										end										
                                    
///////////////////////////////////////////////////////////////////////////////////////////////////////////////         
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
										
									else
										begin
											MoveSpeed = 1 + MoveSpeed_0 + MoveSpeed_1 * 2;
										//Finally getting to the actual tank controls
											if (Up    == 1)
											    begin
												    Tank1_yPos     = Tank1_yPos - MoveSpeed;
												    PrevDirection = Up_Direction;
											    end
											    
											else if (Right == 1)
											    begin
												    Tank1_xPos     = Tank1_xPos + MoveSpeed;
												    PrevDirection = Right_Direction;
											    end
											
											else if (Down  == 1)
											    begin
												    Tank1_yPos     = Tank1_yPos + MoveSpeed;
												    PrevDirection = Down_Direction;		
											    end
											
											else if (Left  == 1)
											    begin
												    Tank1_xPos     = Tank1_xPos - MoveSpeed;  
												    PrevDirection = Left_Direction;		
											    end
										end
								end 	
								
								if(CoinValue[3:0] == 4'b1010) // Get rid of A-F values on segment counter, only display 0-9. 
                                  begin
                                      CoinValue[7:4] = CoinValue[7:4] + 4'b0001;
                                      CoinValue[3:0] = 4'b0000;										      
                                  
                                  end    
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////////////////////////////////         
							xDivPos = ((Val_Row_In[9:5])%20);
                            yDivPos = ((Val_Col_In[9:5])%15);
                            
                            MapArrayData_Y   = MapArray[yDivPos];
                            MapArrayData_X_3 = MapArrayData_Y[4*xDivPos];
                            MapArrayData_X_2 = MapArrayData_Y[4*xDivPos + 1];
                            MapArrayData_X_1 = MapArrayData_Y[4*xDivPos + 2];
                            MapArrayData_X_0 = MapArrayData_Y[4*xDivPos + 3];
                            
                            MapArray_X = {MapArrayData_X_3, MapArrayData_X_2, MapArrayData_X_1, MapArrayData_X_0 };
///////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////// 
                            //within tank bounding box, set image to tank
                            if ((Val_Col_In >= Tank1_yPos) & (Val_Col_In <= Tank1_yPos + TankWidth)
                              & (Val_Row_In >= Tank1_xPos) & (Val_Row_In <= Tank1_xPos + TankWidth))
                                begin
									//If moving upwards, image is normal orientation
									if (PrevDirection == Up_Direction)
										begin
											Tank_XInput = Val_Row_In - Tank1_xPos;
											Tank_YInput = Val_Col_In - Tank1_yPos;
										end
									// If moving downwards, image is mirrored in x
									else if (PrevDirection == Down_Direction)    
										begin
											Tank_XInput = TankWidth - (Val_Row_In - Tank1_xPos)%TankWidth;
											Tank_YInput = TankWidth - (Val_Col_In - Tank1_yPos)%TankWidth;
										end
									// if moving left, image is flipped to horizontal direction
									else if (PrevDirection == Left_Direction)    
										begin
											Tank_YInput = Val_Row_In - Tank1_xPos;
											Tank_XInput = Val_Col_In - Tank1_yPos;
										end
									// if moving right, image is flipped to horizontal, and then mirrored in y 
									else if (PrevDirection == Right_Direction)
										begin
											Tank_YInput = TankWidth - (Val_Row_In - Tank1_xPos)%TankWidth;
											Tank_XInput = TankWidth - (Val_Col_In - Tank1_yPos)%TankWidth;
										end
            
                                    Red   = Colour_Data_Tank[11:8];
                                    Green = Colour_Data_Tank[7:4];
                                    Blue  = Colour_Data_Tank[3:0];
                                
                                end
							//Bullet Draw
							else if (((Val_Col_In >= Bullet_YInput_1 - BulletWidth/2) & (Val_Col_In <= Bullet_YInput_1 + BulletWidth/2))
							       & ((Val_Row_In >= Bullet_XInput_1 - BulletWidth/2) & (Val_Row_In <= Bullet_XInput_1 + BulletWidth/2)))
								begin
								    if (Bullet_Fired_1 == 1)
                                        begin
                                            Red 	= Colour_Data_Bullet[11:8];
                                            Green 	= Colour_Data_Bullet[7:4]; 
                                            Blue 	= Colour_Data_Bullet[3:0]; 
                                        end
                                    else
                                        begin
                                            Red 	= 4'hF;
                                            Green 	= 4'hF;
                                            Blue 	= 4'hF;
                                        end
                                            
								end
							else	
                                //if not within tank bounding box, image is dependant on colour of map.
								//	this will be changed to the colour of specific images dependant on the case	
								//	rather than just flat colours.
                                begin
									case (MapArray_X)
										4'h0:begin  Red   = 4'hF; 
                                                    Green = 4'hF; 
                                                    Blue  = 4'hF; end
										
										4'h1:begin 	Red   = Colour_Data_Solid_Block[11:8];
													Green = Colour_Data_Solid_Block[ 7:4];
													Blue  = Colour_Data_Solid_Block[ 3:0];
										     end
											 
										4'h2:begin  Red   = Colour_Data_Brick[11:8];
													Green = Colour_Data_Brick[ 7:4];
													Blue  = Colour_Data_Brick[ 3:0];
											 end	
											 
										4'h3:begin 
                                                if (ColourSwitch_1 == 0)
                                                    begin
                                                        Red 	= Colour_Data_Coin[11:8];
                                                        Green 	= Colour_Data_Coin[ 7:4];
                                                        Blue 	= Colour_Data_Coin[ 3:0];
                                                    end
                                                else
                                                    begin
                                                        Red 	= Colour_Data_Nyan[11:8];
                                                        Green 	= Colour_Data_Nyan[ 7:4];
                                                        Blue 	= Colour_Data_Nyan[ 3:0];
											         end 
                                            end
										
										4'h4:     begin	Red = 4'hF; Green = 4'h4; Blue = 4'h4; end
										4'h5:     begin	Red = 4'hF; Green = 4'h4; Blue = 4'h4; end
										4'h6:     begin	Red = 4'hF; Green = 4'h4; Blue = 4'h4; end
										4'h7:     begin	Red = 4'hF; Green = 4'h4; Blue = 4'h4; end
										
										default:  begin Red = 4'h8; Green = 4'h8; Blue = 4'h8;end
										
									endcase

            
                                end            
                    end
                
                else
                    begin
                        Red 	= 4'h2;
                        Blue 	= 4'h2;
                        Green 	= 4'h2;
                    end
                end
            end
        end

endmodule
