module Brick_Block(
	input Master_Clock_In,
	input [9 : 0] xInput,
	input [9 : 0] yInput,
	output reg [11:0] ColourData = 12'h000
);

(* rom_style = "block" *)

reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

always @(posedge Master_Clock_In)
	begin


		a = xInput % 32;
		b = yInput % 32;

		Inputs = {a, b};

		case(Inputs)

				20'b000000000000000000 : ColourData = 12'h000;
				20'b000000001000000000 : ColourData = 12'h000;
				20'b000000010000000000 : ColourData = 12'h000;
				20'b000000011000000000 : ColourData = 12'h000;
				20'b000000100000000000 : ColourData = 12'h000;
				20'b000000101000000000 : ColourData = 12'h000;
				20'b000000110000000000 : ColourData = 12'h000;
				20'b000000111000000000 : ColourData = 12'h000;
				20'b000001000000000000 : ColourData = 12'h000;
				20'b000001001000000000 : ColourData = 12'h000;
				20'b000001010000000000 : ColourData = 12'h000;
				20'b000001011000000000 : ColourData = 12'h000;
				20'b000001100000000000 : ColourData = 12'h000;
				20'b000001101000000000 : ColourData = 12'h000;
				20'b000001110000000000 : ColourData = 12'h000;
				20'b000001111000000000 : ColourData = 12'h000;
				20'b000010000000000000 : ColourData = 12'h000;
				20'b000010001000000000 : ColourData = 12'h000;
				20'b000010010000000000 : ColourData = 12'h000;
				20'b000010011000000000 : ColourData = 12'h000;
				20'b000010100000000000 : ColourData = 12'h000;
				20'b000010101000000000 : ColourData = 12'h000;
				20'b000010110000000000 : ColourData = 12'h000;
				20'b000010111000000000 : ColourData = 12'h000;
				20'b000011000000000000 : ColourData = 12'h000;
				20'b000011001000000000 : ColourData = 12'h000;
				20'b000011010000000000 : ColourData = 12'h000;
				20'b000011011000000000 : ColourData = 12'h000;
				20'b000011100000000000 : ColourData = 12'h000;
				20'b000011101000000000 : ColourData = 12'h000;
				20'b000011110000000000 : ColourData = 12'h000;
				20'b000011111000000000 : ColourData = 12'h000;
				20'b000000000000000001 : ColourData = 12'h000;
				20'b000000001000000001 : ColourData = 12'hB75;
				20'b000000010000000001 : ColourData = 12'hB75;
				20'b000000011000000001 : ColourData = 12'hB75;
				20'b000000100000000001 : ColourData = 12'hB75;
				20'b000000101000000001 : ColourData = 12'hB75;
				20'b000000110000000001 : ColourData = 12'hB75;
				20'b000000111000000001 : ColourData = 12'hB75;
				20'b000001000000000001 : ColourData = 12'hB75;
				20'b000001001000000001 : ColourData = 12'hB75;
				20'b000001010000000001 : ColourData = 12'hB75;
				20'b000001011000000001 : ColourData = 12'hB75;
				20'b000001100000000001 : ColourData = 12'hB75;
				20'b000001101000000001 : ColourData = 12'hB75;
				20'b000001110000000001 : ColourData = 12'hB75;
				20'b000001111000000001 : ColourData = 12'h000;
				20'b000010000000000001 : ColourData = 12'h000;
				20'b000010001000000001 : ColourData = 12'hB75;
				20'b000010010000000001 : ColourData = 12'hB75;
				20'b000010011000000001 : ColourData = 12'hB75;
				20'b000010100000000001 : ColourData = 12'hB75;
				20'b000010101000000001 : ColourData = 12'hB75;
				20'b000010110000000001 : ColourData = 12'hB75;
				20'b000010111000000001 : ColourData = 12'hB75;
				20'b000011000000000001 : ColourData = 12'hB75;
				20'b000011001000000001 : ColourData = 12'hB75;
				20'b000011010000000001 : ColourData = 12'hB75;
				20'b000011011000000001 : ColourData = 12'hB75;
				20'b000011100000000001 : ColourData = 12'hB75;
				20'b000011101000000001 : ColourData = 12'hB75;
				20'b000011110000000001 : ColourData = 12'hB75;
				20'b000011111000000001 : ColourData = 12'h000;
				20'b000000000000000010 : ColourData = 12'h000;
				20'b000000001000000010 : ColourData = 12'hB75;
				20'b000000010000000010 : ColourData = 12'h532;
				20'b000000011000000010 : ColourData = 12'h532;
				20'b000000100000000010 : ColourData = 12'h532;
				20'b000000101000000010 : ColourData = 12'h532;
				20'b000000110000000010 : ColourData = 12'h532;
				20'b000000111000000010 : ColourData = 12'h532;
				20'b000001000000000010 : ColourData = 12'h532;
				20'b000001001000000010 : ColourData = 12'h532;
				20'b000001010000000010 : ColourData = 12'h532;
				20'b000001011000000010 : ColourData = 12'h532;
				20'b000001100000000010 : ColourData = 12'h532;
				20'b000001101000000010 : ColourData = 12'h532;
				20'b000001110000000010 : ColourData = 12'h532;
				20'b000001111000000010 : ColourData = 12'h000;
				20'b000010000000000010 : ColourData = 12'h000;
				20'b000010001000000010 : ColourData = 12'hB75;
				20'b000010010000000010 : ColourData = 12'h532;
				20'b000010011000000010 : ColourData = 12'h532;
				20'b000010100000000010 : ColourData = 12'h532;
				20'b000010101000000010 : ColourData = 12'h532;
				20'b000010110000000010 : ColourData = 12'h532;
				20'b000010111000000010 : ColourData = 12'h532;
				20'b000011000000000010 : ColourData = 12'h532;
				20'b000011001000000010 : ColourData = 12'h532;
				20'b000011010000000010 : ColourData = 12'h532;
				20'b000011011000000010 : ColourData = 12'h532;
				20'b000011100000000010 : ColourData = 12'h532;
				20'b000011101000000010 : ColourData = 12'h532;
				20'b000011110000000010 : ColourData = 12'h532;
				20'b000011111000000010 : ColourData = 12'h000;
				20'b000000000000000011 : ColourData = 12'h000;
				20'b000000001000000011 : ColourData = 12'hB75;
				20'b000000010000000011 : ColourData = 12'h532;
				20'b000000011000000011 : ColourData = 12'h532;
				20'b000000100000000011 : ColourData = 12'h532;
				20'b000000101000000011 : ColourData = 12'h532;
				20'b000000110000000011 : ColourData = 12'h532;
				20'b000000111000000011 : ColourData = 12'h532;
				20'b000001000000000011 : ColourData = 12'h532;
				20'b000001001000000011 : ColourData = 12'h532;
				20'b000001010000000011 : ColourData = 12'h532;
				20'b000001011000000011 : ColourData = 12'h532;
				20'b000001100000000011 : ColourData = 12'h532;
				20'b000001101000000011 : ColourData = 12'h532;
				20'b000001110000000011 : ColourData = 12'h532;
				20'b000001111000000011 : ColourData = 12'h000;
				20'b000010000000000011 : ColourData = 12'h000;
				20'b000010001000000011 : ColourData = 12'hB75;
				20'b000010010000000011 : ColourData = 12'h532;
				20'b000010011000000011 : ColourData = 12'h532;
				20'b000010100000000011 : ColourData = 12'h532;
				20'b000010101000000011 : ColourData = 12'h532;
				20'b000010110000000011 : ColourData = 12'h532;
				20'b000010111000000011 : ColourData = 12'h532;
				20'b000011000000000011 : ColourData = 12'h532;
				20'b000011001000000011 : ColourData = 12'h532;
				20'b000011010000000011 : ColourData = 12'h532;
				20'b000011011000000011 : ColourData = 12'h532;
				20'b000011100000000011 : ColourData = 12'h532;
				20'b000011101000000011 : ColourData = 12'h532;
				20'b000011110000000011 : ColourData = 12'h532;
				20'b000011111000000011 : ColourData = 12'h000;
				20'b000000000000000100 : ColourData = 12'h000;
				20'b000000001000000100 : ColourData = 12'hB75;
				20'b000000010000000100 : ColourData = 12'h532;
				20'b000000011000000100 : ColourData = 12'h532;
				20'b000000100000000100 : ColourData = 12'h532;
				20'b000000101000000100 : ColourData = 12'h532;
				20'b000000110000000100 : ColourData = 12'h532;
				20'b000000111000000100 : ColourData = 12'h532;
				20'b000001000000000100 : ColourData = 12'h532;
				20'b000001001000000100 : ColourData = 12'h532;
				20'b000001010000000100 : ColourData = 12'h532;
				20'b000001011000000100 : ColourData = 12'h532;
				20'b000001100000000100 : ColourData = 12'h532;
				20'b000001101000000100 : ColourData = 12'h532;
				20'b000001110000000100 : ColourData = 12'h532;
				20'b000001111000000100 : ColourData = 12'h000;
				20'b000010000000000100 : ColourData = 12'h000;
				20'b000010001000000100 : ColourData = 12'hB75;
				20'b000010010000000100 : ColourData = 12'h532;
				20'b000010011000000100 : ColourData = 12'h532;
				20'b000010100000000100 : ColourData = 12'h532;
				20'b000010101000000100 : ColourData = 12'h532;
				20'b000010110000000100 : ColourData = 12'h532;
				20'b000010111000000100 : ColourData = 12'h532;
				20'b000011000000000100 : ColourData = 12'h532;
				20'b000011001000000100 : ColourData = 12'h532;
				20'b000011010000000100 : ColourData = 12'h532;
				20'b000011011000000100 : ColourData = 12'h532;
				20'b000011100000000100 : ColourData = 12'h532;
				20'b000011101000000100 : ColourData = 12'h532;
				20'b000011110000000100 : ColourData = 12'h532;
				20'b000011111000000100 : ColourData = 12'h000;
				20'b000000000000000101 : ColourData = 12'h000;
				20'b000000001000000101 : ColourData = 12'hB75;
				20'b000000010000000101 : ColourData = 12'h532;
				20'b000000011000000101 : ColourData = 12'h532;
				20'b000000100000000101 : ColourData = 12'h532;
				20'b000000101000000101 : ColourData = 12'h532;
				20'b000000110000000101 : ColourData = 12'h532;
				20'b000000111000000101 : ColourData = 12'h532;
				20'b000001000000000101 : ColourData = 12'h532;
				20'b000001001000000101 : ColourData = 12'h532;
				20'b000001010000000101 : ColourData = 12'h532;
				20'b000001011000000101 : ColourData = 12'h532;
				20'b000001100000000101 : ColourData = 12'h532;
				20'b000001101000000101 : ColourData = 12'h532;
				20'b000001110000000101 : ColourData = 12'h532;
				20'b000001111000000101 : ColourData = 12'h000;
				20'b000010000000000101 : ColourData = 12'h000;
				20'b000010001000000101 : ColourData = 12'hB75;
				20'b000010010000000101 : ColourData = 12'h532;
				20'b000010011000000101 : ColourData = 12'h532;
				20'b000010100000000101 : ColourData = 12'h532;
				20'b000010101000000101 : ColourData = 12'h532;
				20'b000010110000000101 : ColourData = 12'h532;
				20'b000010111000000101 : ColourData = 12'h532;
				20'b000011000000000101 : ColourData = 12'h532;
				20'b000011001000000101 : ColourData = 12'h532;
				20'b000011010000000101 : ColourData = 12'h532;
				20'b000011011000000101 : ColourData = 12'h532;
				20'b000011100000000101 : ColourData = 12'h532;
				20'b000011101000000101 : ColourData = 12'h532;
				20'b000011110000000101 : ColourData = 12'h532;
				20'b000011111000000101 : ColourData = 12'h000;
				20'b000000000000000110 : ColourData = 12'h000;
				20'b000000001000000110 : ColourData = 12'hB75;
				20'b000000010000000110 : ColourData = 12'h532;
				20'b000000011000000110 : ColourData = 12'h532;
				20'b000000100000000110 : ColourData = 12'h532;
				20'b000000101000000110 : ColourData = 12'h532;
				20'b000000110000000110 : ColourData = 12'h532;
				20'b000000111000000110 : ColourData = 12'h532;
				20'b000001000000000110 : ColourData = 12'h532;
				20'b000001001000000110 : ColourData = 12'h532;
				20'b000001010000000110 : ColourData = 12'h532;
				20'b000001011000000110 : ColourData = 12'h532;
				20'b000001100000000110 : ColourData = 12'h532;
				20'b000001101000000110 : ColourData = 12'h532;
				20'b000001110000000110 : ColourData = 12'h532;
				20'b000001111000000110 : ColourData = 12'h000;
				20'b000010000000000110 : ColourData = 12'h000;
				20'b000010001000000110 : ColourData = 12'hB75;
				20'b000010010000000110 : ColourData = 12'h532;
				20'b000010011000000110 : ColourData = 12'h532;
				20'b000010100000000110 : ColourData = 12'h532;
				20'b000010101000000110 : ColourData = 12'h532;
				20'b000010110000000110 : ColourData = 12'h532;
				20'b000010111000000110 : ColourData = 12'h532;
				20'b000011000000000110 : ColourData = 12'h532;
				20'b000011001000000110 : ColourData = 12'h532;
				20'b000011010000000110 : ColourData = 12'h532;
				20'b000011011000000110 : ColourData = 12'h532;
				20'b000011100000000110 : ColourData = 12'h532;
				20'b000011101000000110 : ColourData = 12'h532;
				20'b000011110000000110 : ColourData = 12'h532;
				20'b000011111000000110 : ColourData = 12'h000;
				20'b000000000000000111 : ColourData = 12'h000;
				20'b000000001000000111 : ColourData = 12'h000;
				20'b000000010000000111 : ColourData = 12'h000;
				20'b000000011000000111 : ColourData = 12'h000;
				20'b000000100000000111 : ColourData = 12'h000;
				20'b000000101000000111 : ColourData = 12'h000;
				20'b000000110000000111 : ColourData = 12'h000;
				20'b000000111000000111 : ColourData = 12'h000;
				20'b000001000000000111 : ColourData = 12'h000;
				20'b000001001000000111 : ColourData = 12'h000;
				20'b000001010000000111 : ColourData = 12'h000;
				20'b000001011000000111 : ColourData = 12'h000;
				20'b000001100000000111 : ColourData = 12'h000;
				20'b000001101000000111 : ColourData = 12'h000;
				20'b000001110000000111 : ColourData = 12'h000;
				20'b000001111000000111 : ColourData = 12'h000;
				20'b000010000000000111 : ColourData = 12'h000;
				20'b000010001000000111 : ColourData = 12'h000;
				20'b000010010000000111 : ColourData = 12'h000;
				20'b000010011000000111 : ColourData = 12'h000;
				20'b000010100000000111 : ColourData = 12'h000;
				20'b000010101000000111 : ColourData = 12'h000;
				20'b000010110000000111 : ColourData = 12'h000;
				20'b000010111000000111 : ColourData = 12'h000;
				20'b000011000000000111 : ColourData = 12'h000;
				20'b000011001000000111 : ColourData = 12'h000;
				20'b000011010000000111 : ColourData = 12'h000;
				20'b000011011000000111 : ColourData = 12'h000;
				20'b000011100000000111 : ColourData = 12'h000;
				20'b000011101000000111 : ColourData = 12'h000;
				20'b000011110000000111 : ColourData = 12'h000;
				20'b000011111000000111 : ColourData = 12'h000;
				20'b000000000000001000 : ColourData = 12'h000;
				20'b000000001000001000 : ColourData = 12'h000;
				20'b000000010000001000 : ColourData = 12'h000;
				20'b000000011000001000 : ColourData = 12'h000;
				20'b000000100000001000 : ColourData = 12'h000;
				20'b000000101000001000 : ColourData = 12'h000;
				20'b000000110000001000 : ColourData = 12'h000;
				20'b000000111000001000 : ColourData = 12'h000;
				20'b000001000000001000 : ColourData = 12'h000;
				20'b000001001000001000 : ColourData = 12'h000;
				20'b000001010000001000 : ColourData = 12'h000;
				20'b000001011000001000 : ColourData = 12'h000;
				20'b000001100000001000 : ColourData = 12'h000;
				20'b000001101000001000 : ColourData = 12'h000;
				20'b000001110000001000 : ColourData = 12'h000;
				20'b000001111000001000 : ColourData = 12'h000;
				20'b000010000000001000 : ColourData = 12'h000;
				20'b000010001000001000 : ColourData = 12'h000;
				20'b000010010000001000 : ColourData = 12'h000;
				20'b000010011000001000 : ColourData = 12'h000;
				20'b000010100000001000 : ColourData = 12'h000;
				20'b000010101000001000 : ColourData = 12'h000;
				20'b000010110000001000 : ColourData = 12'h000;
				20'b000010111000001000 : ColourData = 12'h000;
				20'b000011000000001000 : ColourData = 12'h000;
				20'b000011001000001000 : ColourData = 12'h000;
				20'b000011010000001000 : ColourData = 12'h000;
				20'b000011011000001000 : ColourData = 12'h000;
				20'b000011100000001000 : ColourData = 12'h000;
				20'b000011101000001000 : ColourData = 12'h000;
				20'b000011110000001000 : ColourData = 12'h000;
				20'b000011111000001000 : ColourData = 12'h000;
				20'b000000000000001001 : ColourData = 12'hB75;
				20'b000000001000001001 : ColourData = 12'hB75;
				20'b000000010000001001 : ColourData = 12'hB75;
				20'b000000011000001001 : ColourData = 12'hB75;
				20'b000000100000001001 : ColourData = 12'hB75;
				20'b000000101000001001 : ColourData = 12'hB75;
				20'b000000110000001001 : ColourData = 12'hB75;
				20'b000000111000001001 : ColourData = 12'h000;
				20'b000001000000001001 : ColourData = 12'h000;
				20'b000001001000001001 : ColourData = 12'hB75;
				20'b000001010000001001 : ColourData = 12'hB75;
				20'b000001011000001001 : ColourData = 12'hB75;
				20'b000001100000001001 : ColourData = 12'hB75;
				20'b000001101000001001 : ColourData = 12'hB75;
				20'b000001110000001001 : ColourData = 12'hB75;
				20'b000001111000001001 : ColourData = 12'hB75;
				20'b000010000000001001 : ColourData = 12'hB75;
				20'b000010001000001001 : ColourData = 12'hB75;
				20'b000010010000001001 : ColourData = 12'hB75;
				20'b000010011000001001 : ColourData = 12'hB75;
				20'b000010100000001001 : ColourData = 12'hB75;
				20'b000010101000001001 : ColourData = 12'hB75;
				20'b000010110000001001 : ColourData = 12'hB75;
				20'b000010111000001001 : ColourData = 12'h000;
				20'b000011000000001001 : ColourData = 12'h000;
				20'b000011001000001001 : ColourData = 12'hB75;
				20'b000011010000001001 : ColourData = 12'hB75;
				20'b000011011000001001 : ColourData = 12'hB75;
				20'b000011100000001001 : ColourData = 12'hB75;
				20'b000011101000001001 : ColourData = 12'hB75;
				20'b000011110000001001 : ColourData = 12'hB75;
				20'b000011111000001001 : ColourData = 12'hB75;
				20'b000000000000001010 : ColourData = 12'h532;
				20'b000000001000001010 : ColourData = 12'h532;
				20'b000000010000001010 : ColourData = 12'h532;
				20'b000000011000001010 : ColourData = 12'h532;
				20'b000000100000001010 : ColourData = 12'h532;
				20'b000000101000001010 : ColourData = 12'h532;
				20'b000000110000001010 : ColourData = 12'h532;
				20'b000000111000001010 : ColourData = 12'h000;
				20'b000001000000001010 : ColourData = 12'h000;
				20'b000001001000001010 : ColourData = 12'hB75;
				20'b000001010000001010 : ColourData = 12'h532;
				20'b000001011000001010 : ColourData = 12'h532;
				20'b000001100000001010 : ColourData = 12'h532;
				20'b000001101000001010 : ColourData = 12'h532;
				20'b000001110000001010 : ColourData = 12'h532;
				20'b000001111000001010 : ColourData = 12'h532;
				20'b000010000000001010 : ColourData = 12'h532;
				20'b000010001000001010 : ColourData = 12'h532;
				20'b000010010000001010 : ColourData = 12'h532;
				20'b000010011000001010 : ColourData = 12'h532;
				20'b000010100000001010 : ColourData = 12'h532;
				20'b000010101000001010 : ColourData = 12'h532;
				20'b000010110000001010 : ColourData = 12'h532;
				20'b000010111000001010 : ColourData = 12'h000;
				20'b000011000000001010 : ColourData = 12'h000;
				20'b000011001000001010 : ColourData = 12'hB75;
				20'b000011010000001010 : ColourData = 12'h532;
				20'b000011011000001010 : ColourData = 12'h532;
				20'b000011100000001010 : ColourData = 12'h532;
				20'b000011101000001010 : ColourData = 12'h532;
				20'b000011110000001010 : ColourData = 12'h532;
				20'b000011111000001010 : ColourData = 12'h532;
				20'b000000000000001011 : ColourData = 12'h532;
				20'b000000001000001011 : ColourData = 12'h532;
				20'b000000010000001011 : ColourData = 12'h532;
				20'b000000011000001011 : ColourData = 12'h532;
				20'b000000100000001011 : ColourData = 12'h532;
				20'b000000101000001011 : ColourData = 12'h532;
				20'b000000110000001011 : ColourData = 12'h532;
				20'b000000111000001011 : ColourData = 12'h000;
				20'b000001000000001011 : ColourData = 12'h000;
				20'b000001001000001011 : ColourData = 12'hB75;
				20'b000001010000001011 : ColourData = 12'h532;
				20'b000001011000001011 : ColourData = 12'h532;
				20'b000001100000001011 : ColourData = 12'h532;
				20'b000001101000001011 : ColourData = 12'h532;
				20'b000001110000001011 : ColourData = 12'h532;
				20'b000001111000001011 : ColourData = 12'h532;
				20'b000010000000001011 : ColourData = 12'h532;
				20'b000010001000001011 : ColourData = 12'h532;
				20'b000010010000001011 : ColourData = 12'h532;
				20'b000010011000001011 : ColourData = 12'h532;
				20'b000010100000001011 : ColourData = 12'h532;
				20'b000010101000001011 : ColourData = 12'h532;
				20'b000010110000001011 : ColourData = 12'h532;
				20'b000010111000001011 : ColourData = 12'h000;
				20'b000011000000001011 : ColourData = 12'h000;
				20'b000011001000001011 : ColourData = 12'hB75;
				20'b000011010000001011 : ColourData = 12'h532;
				20'b000011011000001011 : ColourData = 12'h532;
				20'b000011100000001011 : ColourData = 12'h532;
				20'b000011101000001011 : ColourData = 12'h532;
				20'b000011110000001011 : ColourData = 12'h532;
				20'b000011111000001011 : ColourData = 12'h532;
				20'b000000000000001100 : ColourData = 12'h532;
				20'b000000001000001100 : ColourData = 12'h532;
				20'b000000010000001100 : ColourData = 12'h532;
				20'b000000011000001100 : ColourData = 12'h532;
				20'b000000100000001100 : ColourData = 12'h532;
				20'b000000101000001100 : ColourData = 12'h532;
				20'b000000110000001100 : ColourData = 12'h532;
				20'b000000111000001100 : ColourData = 12'h000;
				20'b000001000000001100 : ColourData = 12'h000;
				20'b000001001000001100 : ColourData = 12'hB75;
				20'b000001010000001100 : ColourData = 12'h532;
				20'b000001011000001100 : ColourData = 12'h532;
				20'b000001100000001100 : ColourData = 12'h532;
				20'b000001101000001100 : ColourData = 12'h532;
				20'b000001110000001100 : ColourData = 12'h532;
				20'b000001111000001100 : ColourData = 12'h532;
				20'b000010000000001100 : ColourData = 12'h532;
				20'b000010001000001100 : ColourData = 12'h532;
				20'b000010010000001100 : ColourData = 12'h532;
				20'b000010011000001100 : ColourData = 12'h532;
				20'b000010100000001100 : ColourData = 12'h532;
				20'b000010101000001100 : ColourData = 12'h532;
				20'b000010110000001100 : ColourData = 12'h532;
				20'b000010111000001100 : ColourData = 12'h000;
				20'b000011000000001100 : ColourData = 12'h000;
				20'b000011001000001100 : ColourData = 12'hB75;
				20'b000011010000001100 : ColourData = 12'h532;
				20'b000011011000001100 : ColourData = 12'h532;
				20'b000011100000001100 : ColourData = 12'h532;
				20'b000011101000001100 : ColourData = 12'h532;
				20'b000011110000001100 : ColourData = 12'h532;
				20'b000011111000001100 : ColourData = 12'h532;
				20'b000000000000001101 : ColourData = 12'h532;
				20'b000000001000001101 : ColourData = 12'h532;
				20'b000000010000001101 : ColourData = 12'h532;
				20'b000000011000001101 : ColourData = 12'h532;
				20'b000000100000001101 : ColourData = 12'h532;
				20'b000000101000001101 : ColourData = 12'h532;
				20'b000000110000001101 : ColourData = 12'h532;
				20'b000000111000001101 : ColourData = 12'h000;
				20'b000001000000001101 : ColourData = 12'h000;
				20'b000001001000001101 : ColourData = 12'hB75;
				20'b000001010000001101 : ColourData = 12'h532;
				20'b000001011000001101 : ColourData = 12'h532;
				20'b000001100000001101 : ColourData = 12'h532;
				20'b000001101000001101 : ColourData = 12'h532;
				20'b000001110000001101 : ColourData = 12'h532;
				20'b000001111000001101 : ColourData = 12'h532;
				20'b000010000000001101 : ColourData = 12'h532;
				20'b000010001000001101 : ColourData = 12'h532;
				20'b000010010000001101 : ColourData = 12'h532;
				20'b000010011000001101 : ColourData = 12'h532;
				20'b000010100000001101 : ColourData = 12'h532;
				20'b000010101000001101 : ColourData = 12'h532;
				20'b000010110000001101 : ColourData = 12'h532;
				20'b000010111000001101 : ColourData = 12'h000;
				20'b000011000000001101 : ColourData = 12'h000;
				20'b000011001000001101 : ColourData = 12'hB75;
				20'b000011010000001101 : ColourData = 12'h532;
				20'b000011011000001101 : ColourData = 12'h532;
				20'b000011100000001101 : ColourData = 12'h532;
				20'b000011101000001101 : ColourData = 12'h532;
				20'b000011110000001101 : ColourData = 12'h532;
				20'b000011111000001101 : ColourData = 12'h532;
				20'b000000000000001110 : ColourData = 12'h532;
				20'b000000001000001110 : ColourData = 12'h532;
				20'b000000010000001110 : ColourData = 12'h532;
				20'b000000011000001110 : ColourData = 12'h532;
				20'b000000100000001110 : ColourData = 12'h532;
				20'b000000101000001110 : ColourData = 12'h532;
				20'b000000110000001110 : ColourData = 12'h532;
				20'b000000111000001110 : ColourData = 12'h000;
				20'b000001000000001110 : ColourData = 12'h000;
				20'b000001001000001110 : ColourData = 12'hB75;
				20'b000001010000001110 : ColourData = 12'h532;
				20'b000001011000001110 : ColourData = 12'h532;
				20'b000001100000001110 : ColourData = 12'h532;
				20'b000001101000001110 : ColourData = 12'h532;
				20'b000001110000001110 : ColourData = 12'h532;
				20'b000001111000001110 : ColourData = 12'h532;
				20'b000010000000001110 : ColourData = 12'h532;
				20'b000010001000001110 : ColourData = 12'h532;
				20'b000010010000001110 : ColourData = 12'h532;
				20'b000010011000001110 : ColourData = 12'h532;
				20'b000010100000001110 : ColourData = 12'h532;
				20'b000010101000001110 : ColourData = 12'h532;
				20'b000010110000001110 : ColourData = 12'h532;
				20'b000010111000001110 : ColourData = 12'h000;
				20'b000011000000001110 : ColourData = 12'h000;
				20'b000011001000001110 : ColourData = 12'hB75;
				20'b000011010000001110 : ColourData = 12'h532;
				20'b000011011000001110 : ColourData = 12'h532;
				20'b000011100000001110 : ColourData = 12'h532;
				20'b000011101000001110 : ColourData = 12'h532;
				20'b000011110000001110 : ColourData = 12'h532;
				20'b000011111000001110 : ColourData = 12'h532;
				20'b000000000000001111 : ColourData = 12'h000;
				20'b000000001000001111 : ColourData = 12'h000;
				20'b000000010000001111 : ColourData = 12'h000;
				20'b000000011000001111 : ColourData = 12'h000;
				20'b000000100000001111 : ColourData = 12'h000;
				20'b000000101000001111 : ColourData = 12'h000;
				20'b000000110000001111 : ColourData = 12'h000;
				20'b000000111000001111 : ColourData = 12'h000;
				20'b000001000000001111 : ColourData = 12'h000;
				20'b000001001000001111 : ColourData = 12'h000;
				20'b000001010000001111 : ColourData = 12'h000;
				20'b000001011000001111 : ColourData = 12'h000;
				20'b000001100000001111 : ColourData = 12'h000;
				20'b000001101000001111 : ColourData = 12'h000;
				20'b000001110000001111 : ColourData = 12'h000;
				20'b000001111000001111 : ColourData = 12'h000;
				20'b000010000000001111 : ColourData = 12'h000;
				20'b000010001000001111 : ColourData = 12'h000;
				20'b000010010000001111 : ColourData = 12'h000;
				20'b000010011000001111 : ColourData = 12'h000;
				20'b000010100000001111 : ColourData = 12'h000;
				20'b000010101000001111 : ColourData = 12'h000;
				20'b000010110000001111 : ColourData = 12'h000;
				20'b000010111000001111 : ColourData = 12'h000;
				20'b000011000000001111 : ColourData = 12'h000;
				20'b000011001000001111 : ColourData = 12'h000;
				20'b000011010000001111 : ColourData = 12'h000;
				20'b000011011000001111 : ColourData = 12'h000;
				20'b000011100000001111 : ColourData = 12'h000;
				20'b000011101000001111 : ColourData = 12'h000;
				20'b000011110000001111 : ColourData = 12'h000;
				20'b000011111000001111 : ColourData = 12'h000;
				20'b000000000000010000 : ColourData = 12'h000;
				20'b000000001000010000 : ColourData = 12'h000;
				20'b000000010000010000 : ColourData = 12'h000;
				20'b000000011000010000 : ColourData = 12'h000;
				20'b000000100000010000 : ColourData = 12'h000;
				20'b000000101000010000 : ColourData = 12'h000;
				20'b000000110000010000 : ColourData = 12'h000;
				20'b000000111000010000 : ColourData = 12'h000;
				20'b000001000000010000 : ColourData = 12'h000;
				20'b000001001000010000 : ColourData = 12'h000;
				20'b000001010000010000 : ColourData = 12'h000;
				20'b000001011000010000 : ColourData = 12'h000;
				20'b000001100000010000 : ColourData = 12'h000;
				20'b000001101000010000 : ColourData = 12'h000;
				20'b000001110000010000 : ColourData = 12'h000;
				20'b000001111000010000 : ColourData = 12'h000;
				20'b000010000000010000 : ColourData = 12'h000;
				20'b000010001000010000 : ColourData = 12'h000;
				20'b000010010000010000 : ColourData = 12'h000;
				20'b000010011000010000 : ColourData = 12'h000;
				20'b000010100000010000 : ColourData = 12'h000;
				20'b000010101000010000 : ColourData = 12'h000;
				20'b000010110000010000 : ColourData = 12'h000;
				20'b000010111000010000 : ColourData = 12'h000;
				20'b000011000000010000 : ColourData = 12'h000;
				20'b000011001000010000 : ColourData = 12'h000;
				20'b000011010000010000 : ColourData = 12'h000;
				20'b000011011000010000 : ColourData = 12'h000;
				20'b000011100000010000 : ColourData = 12'h000;
				20'b000011101000010000 : ColourData = 12'h000;
				20'b000011110000010000 : ColourData = 12'h000;
				20'b000011111000010000 : ColourData = 12'h000;
				20'b000000000000010001 : ColourData = 12'h000;
				20'b000000001000010001 : ColourData = 12'hB75;
				20'b000000010000010001 : ColourData = 12'hB75;
				20'b000000011000010001 : ColourData = 12'hB75;
				20'b000000100000010001 : ColourData = 12'hB75;
				20'b000000101000010001 : ColourData = 12'hB75;
				20'b000000110000010001 : ColourData = 12'hB75;
				20'b000000111000010001 : ColourData = 12'hB75;
				20'b000001000000010001 : ColourData = 12'hB75;
				20'b000001001000010001 : ColourData = 12'hB75;
				20'b000001010000010001 : ColourData = 12'hB75;
				20'b000001011000010001 : ColourData = 12'hB75;
				20'b000001100000010001 : ColourData = 12'hB75;
				20'b000001101000010001 : ColourData = 12'hB75;
				20'b000001110000010001 : ColourData = 12'hB75;
				20'b000001111000010001 : ColourData = 12'h000;
				20'b000010000000010001 : ColourData = 12'h000;
				20'b000010001000010001 : ColourData = 12'hB75;
				20'b000010010000010001 : ColourData = 12'hB75;
				20'b000010011000010001 : ColourData = 12'hB75;
				20'b000010100000010001 : ColourData = 12'hB75;
				20'b000010101000010001 : ColourData = 12'hB75;
				20'b000010110000010001 : ColourData = 12'hB75;
				20'b000010111000010001 : ColourData = 12'hB75;
				20'b000011000000010001 : ColourData = 12'hB75;
				20'b000011001000010001 : ColourData = 12'hB75;
				20'b000011010000010001 : ColourData = 12'hB75;
				20'b000011011000010001 : ColourData = 12'hB75;
				20'b000011100000010001 : ColourData = 12'hB75;
				20'b000011101000010001 : ColourData = 12'hB75;
				20'b000011110000010001 : ColourData = 12'hB75;
				20'b000011111000010001 : ColourData = 12'h000;
				20'b000000000000010010 : ColourData = 12'h000;
				20'b000000001000010010 : ColourData = 12'hB75;
				20'b000000010000010010 : ColourData = 12'h532;
				20'b000000011000010010 : ColourData = 12'h532;
				20'b000000100000010010 : ColourData = 12'h532;
				20'b000000101000010010 : ColourData = 12'h532;
				20'b000000110000010010 : ColourData = 12'h532;
				20'b000000111000010010 : ColourData = 12'h532;
				20'b000001000000010010 : ColourData = 12'h532;
				20'b000001001000010010 : ColourData = 12'h532;
				20'b000001010000010010 : ColourData = 12'h532;
				20'b000001011000010010 : ColourData = 12'h532;
				20'b000001100000010010 : ColourData = 12'h532;
				20'b000001101000010010 : ColourData = 12'h532;
				20'b000001110000010010 : ColourData = 12'h532;
				20'b000001111000010010 : ColourData = 12'h000;
				20'b000010000000010010 : ColourData = 12'h000;
				20'b000010001000010010 : ColourData = 12'hB75;
				20'b000010010000010010 : ColourData = 12'h532;
				20'b000010011000010010 : ColourData = 12'h532;
				20'b000010100000010010 : ColourData = 12'h532;
				20'b000010101000010010 : ColourData = 12'h532;
				20'b000010110000010010 : ColourData = 12'h532;
				20'b000010111000010010 : ColourData = 12'h532;
				20'b000011000000010010 : ColourData = 12'h532;
				20'b000011001000010010 : ColourData = 12'h532;
				20'b000011010000010010 : ColourData = 12'h532;
				20'b000011011000010010 : ColourData = 12'h532;
				20'b000011100000010010 : ColourData = 12'h532;
				20'b000011101000010010 : ColourData = 12'h532;
				20'b000011110000010010 : ColourData = 12'h532;
				20'b000011111000010010 : ColourData = 12'h000;
				20'b000000000000010011 : ColourData = 12'h000;
				20'b000000001000010011 : ColourData = 12'hB75;
				20'b000000010000010011 : ColourData = 12'h532;
				20'b000000011000010011 : ColourData = 12'h532;
				20'b000000100000010011 : ColourData = 12'h532;
				20'b000000101000010011 : ColourData = 12'h532;
				20'b000000110000010011 : ColourData = 12'h532;
				20'b000000111000010011 : ColourData = 12'h532;
				20'b000001000000010011 : ColourData = 12'h532;
				20'b000001001000010011 : ColourData = 12'h532;
				20'b000001010000010011 : ColourData = 12'h532;
				20'b000001011000010011 : ColourData = 12'h532;
				20'b000001100000010011 : ColourData = 12'h532;
				20'b000001101000010011 : ColourData = 12'h532;
				20'b000001110000010011 : ColourData = 12'h532;
				20'b000001111000010011 : ColourData = 12'h000;
				20'b000010000000010011 : ColourData = 12'h000;
				20'b000010001000010011 : ColourData = 12'hB75;
				20'b000010010000010011 : ColourData = 12'h532;
				20'b000010011000010011 : ColourData = 12'h532;
				20'b000010100000010011 : ColourData = 12'h532;
				20'b000010101000010011 : ColourData = 12'h532;
				20'b000010110000010011 : ColourData = 12'h532;
				20'b000010111000010011 : ColourData = 12'h532;
				20'b000011000000010011 : ColourData = 12'h532;
				20'b000011001000010011 : ColourData = 12'h532;
				20'b000011010000010011 : ColourData = 12'h532;
				20'b000011011000010011 : ColourData = 12'h532;
				20'b000011100000010011 : ColourData = 12'h532;
				20'b000011101000010011 : ColourData = 12'h532;
				20'b000011110000010011 : ColourData = 12'h532;
				20'b000011111000010011 : ColourData = 12'h000;
				20'b000000000000010100 : ColourData = 12'h000;
				20'b000000001000010100 : ColourData = 12'hB75;
				20'b000000010000010100 : ColourData = 12'h532;
				20'b000000011000010100 : ColourData = 12'h532;
				20'b000000100000010100 : ColourData = 12'h532;
				20'b000000101000010100 : ColourData = 12'h532;
				20'b000000110000010100 : ColourData = 12'h532;
				20'b000000111000010100 : ColourData = 12'h532;
				20'b000001000000010100 : ColourData = 12'h532;
				20'b000001001000010100 : ColourData = 12'h532;
				20'b000001010000010100 : ColourData = 12'h532;
				20'b000001011000010100 : ColourData = 12'h532;
				20'b000001100000010100 : ColourData = 12'h532;
				20'b000001101000010100 : ColourData = 12'h532;
				20'b000001110000010100 : ColourData = 12'h532;
				20'b000001111000010100 : ColourData = 12'h000;
				20'b000010000000010100 : ColourData = 12'h000;
				20'b000010001000010100 : ColourData = 12'hB75;
				20'b000010010000010100 : ColourData = 12'h532;
				20'b000010011000010100 : ColourData = 12'h532;
				20'b000010100000010100 : ColourData = 12'h532;
				20'b000010101000010100 : ColourData = 12'h532;
				20'b000010110000010100 : ColourData = 12'h532;
				20'b000010111000010100 : ColourData = 12'h532;
				20'b000011000000010100 : ColourData = 12'h532;
				20'b000011001000010100 : ColourData = 12'h532;
				20'b000011010000010100 : ColourData = 12'h532;
				20'b000011011000010100 : ColourData = 12'h532;
				20'b000011100000010100 : ColourData = 12'h532;
				20'b000011101000010100 : ColourData = 12'h532;
				20'b000011110000010100 : ColourData = 12'h532;
				20'b000011111000010100 : ColourData = 12'h000;
				20'b000000000000010101 : ColourData = 12'h000;
				20'b000000001000010101 : ColourData = 12'hB75;
				20'b000000010000010101 : ColourData = 12'h532;
				20'b000000011000010101 : ColourData = 12'h532;
				20'b000000100000010101 : ColourData = 12'h532;
				20'b000000101000010101 : ColourData = 12'h532;
				20'b000000110000010101 : ColourData = 12'h532;
				20'b000000111000010101 : ColourData = 12'h532;
				20'b000001000000010101 : ColourData = 12'h532;
				20'b000001001000010101 : ColourData = 12'h532;
				20'b000001010000010101 : ColourData = 12'h532;
				20'b000001011000010101 : ColourData = 12'h532;
				20'b000001100000010101 : ColourData = 12'h532;
				20'b000001101000010101 : ColourData = 12'h532;
				20'b000001110000010101 : ColourData = 12'h532;
				20'b000001111000010101 : ColourData = 12'h000;
				20'b000010000000010101 : ColourData = 12'h000;
				20'b000010001000010101 : ColourData = 12'hB75;
				20'b000010010000010101 : ColourData = 12'h532;
				20'b000010011000010101 : ColourData = 12'h532;
				20'b000010100000010101 : ColourData = 12'h532;
				20'b000010101000010101 : ColourData = 12'h532;
				20'b000010110000010101 : ColourData = 12'h532;
				20'b000010111000010101 : ColourData = 12'h532;
				20'b000011000000010101 : ColourData = 12'h532;
				20'b000011001000010101 : ColourData = 12'h532;
				20'b000011010000010101 : ColourData = 12'h532;
				20'b000011011000010101 : ColourData = 12'h532;
				20'b000011100000010101 : ColourData = 12'h532;
				20'b000011101000010101 : ColourData = 12'h532;
				20'b000011110000010101 : ColourData = 12'h532;
				20'b000011111000010101 : ColourData = 12'h000;
				20'b000000000000010110 : ColourData = 12'h000;
				20'b000000001000010110 : ColourData = 12'hB75;
				20'b000000010000010110 : ColourData = 12'h532;
				20'b000000011000010110 : ColourData = 12'h532;
				20'b000000100000010110 : ColourData = 12'h532;
				20'b000000101000010110 : ColourData = 12'h532;
				20'b000000110000010110 : ColourData = 12'h532;
				20'b000000111000010110 : ColourData = 12'h532;
				20'b000001000000010110 : ColourData = 12'h532;
				20'b000001001000010110 : ColourData = 12'h532;
				20'b000001010000010110 : ColourData = 12'h532;
				20'b000001011000010110 : ColourData = 12'h532;
				20'b000001100000010110 : ColourData = 12'h532;
				20'b000001101000010110 : ColourData = 12'h532;
				20'b000001110000010110 : ColourData = 12'h532;
				20'b000001111000010110 : ColourData = 12'h000;
				20'b000010000000010110 : ColourData = 12'h000;
				20'b000010001000010110 : ColourData = 12'hB75;
				20'b000010010000010110 : ColourData = 12'h532;
				20'b000010011000010110 : ColourData = 12'h532;
				20'b000010100000010110 : ColourData = 12'h532;
				20'b000010101000010110 : ColourData = 12'h532;
				20'b000010110000010110 : ColourData = 12'h532;
				20'b000010111000010110 : ColourData = 12'h532;
				20'b000011000000010110 : ColourData = 12'h532;
				20'b000011001000010110 : ColourData = 12'h532;
				20'b000011010000010110 : ColourData = 12'h532;
				20'b000011011000010110 : ColourData = 12'h532;
				20'b000011100000010110 : ColourData = 12'h532;
				20'b000011101000010110 : ColourData = 12'h532;
				20'b000011110000010110 : ColourData = 12'h532;
				20'b000011111000010110 : ColourData = 12'h000;
				20'b000000000000010111 : ColourData = 12'h000;
				20'b000000001000010111 : ColourData = 12'h000;
				20'b000000010000010111 : ColourData = 12'h000;
				20'b000000011000010111 : ColourData = 12'h000;
				20'b000000100000010111 : ColourData = 12'h000;
				20'b000000101000010111 : ColourData = 12'h000;
				20'b000000110000010111 : ColourData = 12'h000;
				20'b000000111000010111 : ColourData = 12'h000;
				20'b000001000000010111 : ColourData = 12'h000;
				20'b000001001000010111 : ColourData = 12'h000;
				20'b000001010000010111 : ColourData = 12'h000;
				20'b000001011000010111 : ColourData = 12'h000;
				20'b000001100000010111 : ColourData = 12'h000;
				20'b000001101000010111 : ColourData = 12'h000;
				20'b000001110000010111 : ColourData = 12'h000;
				20'b000001111000010111 : ColourData = 12'h000;
				20'b000010000000010111 : ColourData = 12'h000;
				20'b000010001000010111 : ColourData = 12'h000;
				20'b000010010000010111 : ColourData = 12'h000;
				20'b000010011000010111 : ColourData = 12'h000;
				20'b000010100000010111 : ColourData = 12'h000;
				20'b000010101000010111 : ColourData = 12'h000;
				20'b000010110000010111 : ColourData = 12'h000;
				20'b000010111000010111 : ColourData = 12'h000;
				20'b000011000000010111 : ColourData = 12'h000;
				20'b000011001000010111 : ColourData = 12'h000;
				20'b000011010000010111 : ColourData = 12'h000;
				20'b000011011000010111 : ColourData = 12'h000;
				20'b000011100000010111 : ColourData = 12'h000;
				20'b000011101000010111 : ColourData = 12'h000;
				20'b000011110000010111 : ColourData = 12'h000;
				20'b000011111000010111 : ColourData = 12'h000;
				20'b000000000000011000 : ColourData = 12'h000;
				20'b000000001000011000 : ColourData = 12'h000;
				20'b000000010000011000 : ColourData = 12'h000;
				20'b000000011000011000 : ColourData = 12'h000;
				20'b000000100000011000 : ColourData = 12'h000;
				20'b000000101000011000 : ColourData = 12'h000;
				20'b000000110000011000 : ColourData = 12'h000;
				20'b000000111000011000 : ColourData = 12'h000;
				20'b000001000000011000 : ColourData = 12'h000;
				20'b000001001000011000 : ColourData = 12'h000;
				20'b000001010000011000 : ColourData = 12'h000;
				20'b000001011000011000 : ColourData = 12'h000;
				20'b000001100000011000 : ColourData = 12'h000;
				20'b000001101000011000 : ColourData = 12'h000;
				20'b000001110000011000 : ColourData = 12'h000;
				20'b000001111000011000 : ColourData = 12'h000;
				20'b000010000000011000 : ColourData = 12'h000;
				20'b000010001000011000 : ColourData = 12'h000;
				20'b000010010000011000 : ColourData = 12'h000;
				20'b000010011000011000 : ColourData = 12'h000;
				20'b000010100000011000 : ColourData = 12'h000;
				20'b000010101000011000 : ColourData = 12'h000;
				20'b000010110000011000 : ColourData = 12'h000;
				20'b000010111000011000 : ColourData = 12'h000;
				20'b000011000000011000 : ColourData = 12'h000;
				20'b000011001000011000 : ColourData = 12'h000;
				20'b000011010000011000 : ColourData = 12'h000;
				20'b000011011000011000 : ColourData = 12'h000;
				20'b000011100000011000 : ColourData = 12'h000;
				20'b000011101000011000 : ColourData = 12'h000;
				20'b000011110000011000 : ColourData = 12'h000;
				20'b000011111000011000 : ColourData = 12'h000;
				20'b000000000000011001 : ColourData = 12'hB75;
				20'b000000001000011001 : ColourData = 12'hB75;
				20'b000000010000011001 : ColourData = 12'hB75;
				20'b000000011000011001 : ColourData = 12'hB75;
				20'b000000100000011001 : ColourData = 12'hB75;
				20'b000000101000011001 : ColourData = 12'hB75;
				20'b000000110000011001 : ColourData = 12'hB75;
				20'b000000111000011001 : ColourData = 12'h000;
				20'b000001000000011001 : ColourData = 12'h000;
				20'b000001001000011001 : ColourData = 12'hB75;
				20'b000001010000011001 : ColourData = 12'hB75;
				20'b000001011000011001 : ColourData = 12'hB75;
				20'b000001100000011001 : ColourData = 12'hB75;
				20'b000001101000011001 : ColourData = 12'hB75;
				20'b000001110000011001 : ColourData = 12'hB75;
				20'b000001111000011001 : ColourData = 12'hB75;
				20'b000010000000011001 : ColourData = 12'hB75;
				20'b000010001000011001 : ColourData = 12'hB75;
				20'b000010010000011001 : ColourData = 12'hB75;
				20'b000010011000011001 : ColourData = 12'hB75;
				20'b000010100000011001 : ColourData = 12'hB75;
				20'b000010101000011001 : ColourData = 12'hB75;
				20'b000010110000011001 : ColourData = 12'hB75;
				20'b000010111000011001 : ColourData = 12'h000;
				20'b000011000000011001 : ColourData = 12'h000;
				20'b000011001000011001 : ColourData = 12'hB75;
				20'b000011010000011001 : ColourData = 12'hB75;
				20'b000011011000011001 : ColourData = 12'hB75;
				20'b000011100000011001 : ColourData = 12'hB75;
				20'b000011101000011001 : ColourData = 12'hB75;
				20'b000011110000011001 : ColourData = 12'hB75;
				20'b000011111000011001 : ColourData = 12'hB75;
				20'b000000000000011010 : ColourData = 12'h532;
				20'b000000001000011010 : ColourData = 12'h532;
				20'b000000010000011010 : ColourData = 12'h532;
				20'b000000011000011010 : ColourData = 12'h532;
				20'b000000100000011010 : ColourData = 12'h532;
				20'b000000101000011010 : ColourData = 12'h532;
				20'b000000110000011010 : ColourData = 12'h532;
				20'b000000111000011010 : ColourData = 12'h000;
				20'b000001000000011010 : ColourData = 12'h000;
				20'b000001001000011010 : ColourData = 12'hB75;
				20'b000001010000011010 : ColourData = 12'h532;
				20'b000001011000011010 : ColourData = 12'h532;
				20'b000001100000011010 : ColourData = 12'h532;
				20'b000001101000011010 : ColourData = 12'h532;
				20'b000001110000011010 : ColourData = 12'h532;
				20'b000001111000011010 : ColourData = 12'h532;
				20'b000010000000011010 : ColourData = 12'h532;
				20'b000010001000011010 : ColourData = 12'h532;
				20'b000010010000011010 : ColourData = 12'h532;
				20'b000010011000011010 : ColourData = 12'h532;
				20'b000010100000011010 : ColourData = 12'h532;
				20'b000010101000011010 : ColourData = 12'h532;
				20'b000010110000011010 : ColourData = 12'h532;
				20'b000010111000011010 : ColourData = 12'h000;
				20'b000011000000011010 : ColourData = 12'h000;
				20'b000011001000011010 : ColourData = 12'hB75;
				20'b000011010000011010 : ColourData = 12'h532;
				20'b000011011000011010 : ColourData = 12'h532;
				20'b000011100000011010 : ColourData = 12'h532;
				20'b000011101000011010 : ColourData = 12'h532;
				20'b000011110000011010 : ColourData = 12'h532;
				20'b000011111000011010 : ColourData = 12'h532;
				20'b000000000000011011 : ColourData = 12'h532;
				20'b000000001000011011 : ColourData = 12'h532;
				20'b000000010000011011 : ColourData = 12'h532;
				20'b000000011000011011 : ColourData = 12'h532;
				20'b000000100000011011 : ColourData = 12'h532;
				20'b000000101000011011 : ColourData = 12'h532;
				20'b000000110000011011 : ColourData = 12'h532;
				20'b000000111000011011 : ColourData = 12'h000;
				20'b000001000000011011 : ColourData = 12'h000;
				20'b000001001000011011 : ColourData = 12'hB75;
				20'b000001010000011011 : ColourData = 12'h532;
				20'b000001011000011011 : ColourData = 12'h532;
				20'b000001100000011011 : ColourData = 12'h532;
				20'b000001101000011011 : ColourData = 12'h532;
				20'b000001110000011011 : ColourData = 12'h532;
				20'b000001111000011011 : ColourData = 12'h532;
				20'b000010000000011011 : ColourData = 12'h532;
				20'b000010001000011011 : ColourData = 12'h532;
				20'b000010010000011011 : ColourData = 12'h532;
				20'b000010011000011011 : ColourData = 12'h532;
				20'b000010100000011011 : ColourData = 12'h532;
				20'b000010101000011011 : ColourData = 12'h532;
				20'b000010110000011011 : ColourData = 12'h532;
				20'b000010111000011011 : ColourData = 12'h000;
				20'b000011000000011011 : ColourData = 12'h000;
				20'b000011001000011011 : ColourData = 12'hB75;
				20'b000011010000011011 : ColourData = 12'h532;
				20'b000011011000011011 : ColourData = 12'h532;
				20'b000011100000011011 : ColourData = 12'h532;
				20'b000011101000011011 : ColourData = 12'h532;
				20'b000011110000011011 : ColourData = 12'h532;
				20'b000011111000011011 : ColourData = 12'h532;
				20'b000000000000011100 : ColourData = 12'h532;
				20'b000000001000011100 : ColourData = 12'h532;
				20'b000000010000011100 : ColourData = 12'h532;
				20'b000000011000011100 : ColourData = 12'h532;
				20'b000000100000011100 : ColourData = 12'h532;
				20'b000000101000011100 : ColourData = 12'h532;
				20'b000000110000011100 : ColourData = 12'h532;
				20'b000000111000011100 : ColourData = 12'h000;
				20'b000001000000011100 : ColourData = 12'h000;
				20'b000001001000011100 : ColourData = 12'hB75;
				20'b000001010000011100 : ColourData = 12'h532;
				20'b000001011000011100 : ColourData = 12'h532;
				20'b000001100000011100 : ColourData = 12'h532;
				20'b000001101000011100 : ColourData = 12'h532;
				20'b000001110000011100 : ColourData = 12'h532;
				20'b000001111000011100 : ColourData = 12'h532;
				20'b000010000000011100 : ColourData = 12'h532;
				20'b000010001000011100 : ColourData = 12'h532;
				20'b000010010000011100 : ColourData = 12'h532;
				20'b000010011000011100 : ColourData = 12'h532;
				20'b000010100000011100 : ColourData = 12'h532;
				20'b000010101000011100 : ColourData = 12'h532;
				20'b000010110000011100 : ColourData = 12'h532;
				20'b000010111000011100 : ColourData = 12'h000;
				20'b000011000000011100 : ColourData = 12'h000;
				20'b000011001000011100 : ColourData = 12'hB75;
				20'b000011010000011100 : ColourData = 12'h532;
				20'b000011011000011100 : ColourData = 12'h532;
				20'b000011100000011100 : ColourData = 12'h532;
				20'b000011101000011100 : ColourData = 12'h532;
				20'b000011110000011100 : ColourData = 12'h532;
				20'b000011111000011100 : ColourData = 12'h532;
				20'b000000000000011101 : ColourData = 12'h532;
				20'b000000001000011101 : ColourData = 12'h532;
				20'b000000010000011101 : ColourData = 12'h532;
				20'b000000011000011101 : ColourData = 12'h532;
				20'b000000100000011101 : ColourData = 12'h532;
				20'b000000101000011101 : ColourData = 12'h532;
				20'b000000110000011101 : ColourData = 12'h532;
				20'b000000111000011101 : ColourData = 12'h000;
				20'b000001000000011101 : ColourData = 12'h000;
				20'b000001001000011101 : ColourData = 12'hB75;
				20'b000001010000011101 : ColourData = 12'h532;
				20'b000001011000011101 : ColourData = 12'h532;
				20'b000001100000011101 : ColourData = 12'h532;
				20'b000001101000011101 : ColourData = 12'h532;
				20'b000001110000011101 : ColourData = 12'h532;
				20'b000001111000011101 : ColourData = 12'h532;
				20'b000010000000011101 : ColourData = 12'h532;
				20'b000010001000011101 : ColourData = 12'h532;
				20'b000010010000011101 : ColourData = 12'h532;
				20'b000010011000011101 : ColourData = 12'h532;
				20'b000010100000011101 : ColourData = 12'h532;
				20'b000010101000011101 : ColourData = 12'h532;
				20'b000010110000011101 : ColourData = 12'h532;
				20'b000010111000011101 : ColourData = 12'h000;
				20'b000011000000011101 : ColourData = 12'h000;
				20'b000011001000011101 : ColourData = 12'hB75;
				20'b000011010000011101 : ColourData = 12'h532;
				20'b000011011000011101 : ColourData = 12'h532;
				20'b000011100000011101 : ColourData = 12'h532;
				20'b000011101000011101 : ColourData = 12'h532;
				20'b000011110000011101 : ColourData = 12'h532;
				20'b000011111000011101 : ColourData = 12'h532;
				20'b000000000000011110 : ColourData = 12'h532;
				20'b000000001000011110 : ColourData = 12'h532;
				20'b000000010000011110 : ColourData = 12'h532;
				20'b000000011000011110 : ColourData = 12'h532;
				20'b000000100000011110 : ColourData = 12'h532;
				20'b000000101000011110 : ColourData = 12'h532;
				20'b000000110000011110 : ColourData = 12'h532;
				20'b000000111000011110 : ColourData = 12'h000;
				20'b000001000000011110 : ColourData = 12'h000;
				20'b000001001000011110 : ColourData = 12'hB75;
				20'b000001010000011110 : ColourData = 12'h532;
				20'b000001011000011110 : ColourData = 12'h532;
				20'b000001100000011110 : ColourData = 12'h532;
				20'b000001101000011110 : ColourData = 12'h532;
				20'b000001110000011110 : ColourData = 12'h532;
				20'b000001111000011110 : ColourData = 12'h532;
				20'b000010000000011110 : ColourData = 12'h532;
				20'b000010001000011110 : ColourData = 12'h532;
				20'b000010010000011110 : ColourData = 12'h532;
				20'b000010011000011110 : ColourData = 12'h532;
				20'b000010100000011110 : ColourData = 12'h532;
				20'b000010101000011110 : ColourData = 12'h532;
				20'b000010110000011110 : ColourData = 12'h532;
				20'b000010111000011110 : ColourData = 12'h000;
				20'b000011000000011110 : ColourData = 12'h000;
				20'b000011001000011110 : ColourData = 12'hB75;
				20'b000011010000011110 : ColourData = 12'h532;
				20'b000011011000011110 : ColourData = 12'h532;
				20'b000011100000011110 : ColourData = 12'h532;
				20'b000011101000011110 : ColourData = 12'h532;
				20'b000011110000011110 : ColourData = 12'h532;
				20'b000011111000011110 : ColourData = 12'h532;
				20'b000000000000011111 : ColourData = 12'h000;
				20'b000000001000011111 : ColourData = 12'h000;
				20'b000000010000011111 : ColourData = 12'h000;
				20'b000000011000011111 : ColourData = 12'h000;
				20'b000000100000011111 : ColourData = 12'h000;
				20'b000000101000011111 : ColourData = 12'h000;
				20'b000000110000011111 : ColourData = 12'h000;
				20'b000000111000011111 : ColourData = 12'h000;
				20'b000001000000011111 : ColourData = 12'h000;
				20'b000001001000011111 : ColourData = 12'h000;
				20'b000001010000011111 : ColourData = 12'h000;
				20'b000001011000011111 : ColourData = 12'h000;
				20'b000001100000011111 : ColourData = 12'h000;
				20'b000001101000011111 : ColourData = 12'h000;
				20'b000001110000011111 : ColourData = 12'h000;
				20'b000001111000011111 : ColourData = 12'h000;
				20'b000010000000011111 : ColourData = 12'h000;
				20'b000010001000011111 : ColourData = 12'h000;
				20'b000010010000011111 : ColourData = 12'h000;
				20'b000010011000011111 : ColourData = 12'h000;
				20'b000010100000011111 : ColourData = 12'h000;
				20'b000010101000011111 : ColourData = 12'h000;
				20'b000010110000011111 : ColourData = 12'h000;
				20'b000010111000011111 : ColourData = 12'h000;
				20'b000011000000011111 : ColourData = 12'h000;
				20'b000011001000011111 : ColourData = 12'h000;
				20'b000011010000011111 : ColourData = 12'h000;
				20'b000011011000011111 : ColourData = 12'h000;
				20'b000011100000011111 : ColourData = 12'h000;
				20'b000011101000011111 : ColourData = 12'h000;
				20'b000011110000011111 : ColourData = 12'h000;
				20'b000011111000011111 : ColourData = 12'h000;

			endcase		
		end

endmodule

