
//////////////////////////////////////////////////////////////////////////////////
//Map file for bullet
//////////////////////////////////////////////////////////////////////////////////


module Bullet(

  input Master_Clock_In,
  input [9 : 0] xInput,
  input [9 : 0] yInput,
  output reg [11:0] ColourData = 12'h000

);

(* rom_style = "block" *)

reg [19:0] Inputs = 20'd0;

reg [9:0] a, b = 10'd0;

always @(posedge Master_Clock_In)
begin
  a = xInput % 10;
  b = yInput % 10;

Inputs = {a, b};

    case(Inputs)    


20'b00000000000000000000 : ColourData = 12'hFFF;
20'b00000000010000000000 : ColourData = 12'hFFF;
20'b00000000100000000000 : ColourData = 12'h222;
20'b00000000110000000000 : ColourData = 12'h222;
20'b00000001000000000000 : ColourData = 12'h222;
20'b00000001010000000000 : ColourData = 12'h222;
20'b00000001100000000000 : ColourData = 12'h222;
20'b00000001110000000000 : ColourData = 12'h222;
20'b00000010000000000000 : ColourData = 12'hFFF;
20'b00000010010000000000 : ColourData = 12'hFFF;
20'b00000000000000000001 : ColourData = 12'hFFF;
20'b00000000010000000001 : ColourData = 12'h222;
20'b00000000100000000001 : ColourData = 12'h222;
20'b00000000110000000001 : ColourData = 12'h222;
20'b00000001000000000001 : ColourData = 12'h222;
20'b00000001010000000001 : ColourData = 12'h222;
20'b00000001100000000001 : ColourData = 12'h222;
20'b00000001110000000001 : ColourData = 12'h222;
20'b00000010000000000001 : ColourData = 12'h222;
20'b00000010010000000001 : ColourData = 12'hFFF;
20'b00000000000000000010 : ColourData = 12'h222;
20'b00000000010000000010 : ColourData = 12'h222;
20'b00000000100000000010 : ColourData = 12'h222;
20'b00000000110000000010 : ColourData = 12'h222;
20'b00000001000000000010 : ColourData = 12'h000;
20'b00000001010000000010 : ColourData = 12'h000;
20'b00000001100000000010 : ColourData = 12'h222;
20'b00000001110000000010 : ColourData = 12'h222;
20'b00000010000000000010 : ColourData = 12'h222;
20'b00000010010000000010 : ColourData = 12'h222;
20'b00000000000000000011 : ColourData = 12'h222;
20'b00000000010000000011 : ColourData = 12'h222;
20'b00000000100000000011 : ColourData = 12'h222;
20'b00000000110000000011 : ColourData = 12'h000;
20'b00000001000000000011 : ColourData = 12'h000;
20'b00000001010000000011 : ColourData = 12'h000;
20'b00000001100000000011 : ColourData = 12'h000;
20'b00000001110000000011 : ColourData = 12'h222;
20'b00000010000000000011 : ColourData = 12'h222;
20'b00000010010000000011 : ColourData = 12'h222;
20'b00000000000000000100 : ColourData = 12'h222;
20'b00000000010000000100 : ColourData = 12'h222;
20'b00000000100000000100 : ColourData = 12'h000;
20'b00000000110000000100 : ColourData = 12'h000;
20'b00000001000000000100 : ColourData = 12'hFFF;
20'b00000001010000000100 : ColourData = 12'h000;
20'b00000001100000000100 : ColourData = 12'h000;
20'b00000001110000000100 : ColourData = 12'h000;
20'b00000010000000000100 : ColourData = 12'h222;
20'b00000010010000000100 : ColourData = 12'h222;
20'b00000000000000000101 : ColourData = 12'h222;
20'b00000000010000000101 : ColourData = 12'h222;
20'b00000000100000000101 : ColourData = 12'h000;
20'b00000000110000000101 : ColourData = 12'h000;
20'b00000001000000000101 : ColourData = 12'h000;
20'b00000001010000000101 : ColourData = 12'h000;
20'b00000001100000000101 : ColourData = 12'h000;
20'b00000001110000000101 : ColourData = 12'h000;
20'b00000010000000000101 : ColourData = 12'h222;
20'b00000010010000000101 : ColourData = 12'h222;
20'b00000000000000000110 : ColourData = 12'h222;
20'b00000000010000000110 : ColourData = 12'h222;
20'b00000000100000000110 : ColourData = 12'h222;
20'b00000000110000000110 : ColourData = 12'h000;
20'b00000001000000000110 : ColourData = 12'h000;
20'b00000001010000000110 : ColourData = 12'h000;
20'b00000001100000000110 : ColourData = 12'h000;
20'b00000001110000000110 : ColourData = 12'h222;
20'b00000010000000000110 : ColourData = 12'h222;
20'b00000010010000000110 : ColourData = 12'h222;
20'b00000000000000000111 : ColourData = 12'h222;
20'b00000000010000000111 : ColourData = 12'h222;
20'b00000000100000000111 : ColourData = 12'h222;
20'b00000000110000000111 : ColourData = 12'h222;
20'b00000001000000000111 : ColourData = 12'h000;
20'b00000001010000000111 : ColourData = 12'h000;
20'b00000001100000000111 : ColourData = 12'h222;
20'b00000001110000000111 : ColourData = 12'h222;
20'b00000010000000000111 : ColourData = 12'h222;
20'b00000010010000000111 : ColourData = 12'h222;
20'b00000000000000001000 : ColourData = 12'hFFF;
20'b00000000010000001000 : ColourData = 12'h222;
20'b00000000100000001000 : ColourData = 12'h222;
20'b00000000110000001000 : ColourData = 12'h222;
20'b00000001000000001000 : ColourData = 12'h222;
20'b00000001010000001000 : ColourData = 12'h222;
20'b00000001100000001000 : ColourData = 12'h222;
20'b00000001110000001000 : ColourData = 12'h222;
20'b00000010000000001000 : ColourData = 12'h222;
20'b00000010010000001000 : ColourData = 12'hFFF;
20'b00000000000000001001 : ColourData = 12'hFFF;
20'b00000000010000001001 : ColourData = 12'hFFF;
20'b00000000100000001001 : ColourData = 12'h222;
20'b00000000110000001001 : ColourData = 12'h222;
20'b00000001000000001001 : ColourData = 12'h222;
20'b00000001010000001001 : ColourData = 12'h222;
20'b00000001100000001001 : ColourData = 12'h222;
20'b00000001110000001001 : ColourData = 12'h222;
20'b00000010000000001001 : ColourData = 12'hFFF;
20'b00000010010000001001 : ColourData = 12'hFFF;


default: ColourData = 12'h000;

endcase
end

endmodule
